parameter integer matrixH [0:10757] = {
/* num inputs = 360(in0-in359) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 25 */
//* total number of input in adders 3425 */

/* out0000_em-eta0-phi0*/	0,
/* out0001_em-eta1-phi0*/	0,
/* out0002_em-eta2-phi0*/	0,
/* out0003_em-eta3-phi0*/	0,
/* out0004_em-eta4-phi0*/	3,238,0,7,238,1,1,268,2,2,
/* out0005_em-eta5-phi0*/	4,238,0,9,238,1,14,238,2,9,268,2,1,
/* out0006_em-eta6-phi0*/	6,206,0,16,206,1,9,206,2,2,238,2,7,242,0,1,242,2,1,
/* out0007_em-eta7-phi0*/	4,172,0,11,172,1,1,206,1,3,206,2,14,
/* out0008_em-eta8-phi0*/	3,172,0,5,172,1,6,172,2,8,
/* out0009_em-eta9-phi0*/	3,140,0,10,140,1,1,172,2,5,
/* out0010_em-eta10-phi0*/	4,140,0,3,140,1,3,140,2,8,264,0,1,
/* out0011_em-eta11-phi0*/	7,106,0,7,140,2,4,228,4,15,228,5,2,229,0,5,229,1,16,264,0,3,
/* out0012_em-eta12-phi0*/	11,84,4,15,85,0,3,85,1,4,120,0,4,106,0,5,106,1,1,106,2,4,228,5,6,229,0,11,229,4,8,229,5,3,
/* out0013_em-eta13-phi0*/	11,74,0,1,106,2,7,84,5,8,85,0,13,85,1,12,85,4,10,85,5,2,229,2,12,229,3,4,229,4,8,229,5,4,
/* out0014_em-eta14-phi0*/	13,74,0,7,85,2,10,85,3,4,85,4,6,85,5,4,192,4,12,192,5,1,193,0,1,193,1,16,229,2,2,229,3,12,336,4,3,337,1,12,
/* out0015_em-eta15-phi0*/	14,48,4,12,49,1,4,85,2,4,85,3,12,74,0,2,74,2,4,192,5,3,193,0,12,193,4,3,336,4,9,336,5,2,337,0,4,337,1,4,352,0,4,
/* out0016_em-eta16-phi0*/	13,48,5,3,49,0,12,49,1,12,49,4,1,74,2,5,193,2,1,193,3,13,193,4,10,193,5,2,336,5,1,337,0,9,337,4,6,352,0,5,
/* out0017_em-eta17-phi0*/	14,44,2,5,74,2,1,49,2,1,49,3,1,49,4,11,49,5,2,163,3,2,193,2,8,193,3,3,337,2,3,337,3,3,337,4,6,337,5,2,352,0,2,
/* out0018_em-eta18-phi0*/	13,19,3,2,49,2,8,49,3,4,44,0,1,44,2,3,162,2,10,162,3,4,163,3,12,163,4,4,307,3,10,337,2,6,337,3,13,334,2,2,
/* out0019_em-eta19-phi0*/	19,18,2,16,18,3,4,19,3,12,19,4,16,49,3,11,44,0,1,162,0,5,162,1,16,162,2,6,162,3,1,163,4,12,306,0,1,306,1,16,306,2,16,306,3,5,307,3,5,307,4,16,334,0,1,334,2,2,
/* out0020_em-eta0-phi1*/	0,
/* out0021_em-eta1-phi1*/	0,
/* out0022_em-eta2-phi1*/	0,
/* out0023_em-eta3-phi1*/	0,
/* out0024_em-eta4-phi1*/	2,268,1,3,268,2,8,
/* out0025_em-eta5-phi1*/	5,238,1,1,242,0,14,242,1,4,268,1,11,268,2,5,
/* out0026_em-eta6-phi1*/	5,206,1,3,208,0,5,242,0,1,242,1,2,242,2,15,
/* out0027_em-eta7-phi1*/	5,172,1,1,206,1,1,208,0,10,208,1,1,208,2,9,
/* out0028_em-eta8-phi1*/	3,172,1,7,176,0,8,208,2,4,
/* out0029_em-eta9-phi1*/	7,140,0,3,140,1,4,172,1,1,172,2,3,176,0,3,176,2,8,265,1,1,
/* out0030_em-eta10-phi1*/	9,140,1,8,140,2,3,142,0,4,176,2,1,264,0,3,264,1,15,264,2,5,265,0,2,265,1,11,
/* out0031_em-eta11-phi1*/	17,106,0,4,106,1,3,140,2,1,142,0,2,142,2,3,120,0,2,120,1,14,120,2,3,121,0,2,121,1,12,228,4,1,228,5,1,264,0,9,264,1,1,264,2,9,264,3,12,265,3,1,
/* out0032_em-eta12-phi1*/	14,84,4,1,120,0,10,120,1,2,120,2,11,120,3,10,121,3,1,106,1,9,106,2,2,228,5,7,229,5,7,234,1,4,235,1,2,264,3,4,265,3,3,
/* out0033_em-eta13-phi1*/	16,74,0,1,106,1,2,106,2,3,110,0,1,110,2,1,84,5,8,85,5,6,90,1,3,91,1,3,120,3,6,121,3,4,229,2,2,229,5,2,234,0,8,234,1,10,234,2,1,
/* out0034_em-eta14-phi1*/	11,74,0,4,74,1,4,85,2,2,85,5,4,90,0,6,90,1,11,192,4,4,192,5,1,234,0,8,234,3,6,352,1,1,
/* out0035_em-eta15-phi1*/	16,48,4,4,90,0,10,90,2,1,90,3,5,74,0,1,74,1,5,74,2,1,192,5,11,193,0,3,193,4,1,193,5,4,234,3,1,336,4,4,336,5,5,352,0,1,352,1,7,
/* out0036_em-eta16-phi1*/	20,44,2,1,74,1,1,74,2,4,48,5,12,49,0,4,49,4,1,49,5,2,90,3,2,193,2,2,193,4,2,193,5,9,198,0,1,198,1,1,336,5,8,337,0,3,337,4,4,337,5,7,352,0,3,352,1,1,352,2,3,
/* out0037_em-eta17-phi1*/	17,44,0,1,44,2,4,74,2,1,49,2,1,49,4,3,49,5,11,54,1,1,163,3,1,193,2,5,198,0,6,334,2,1,352,0,1,352,2,4,337,2,4,337,5,6,342,0,2,342,1,1,
/* out0038_em-eta18-phi1*/	15,18,3,1,19,3,1,49,2,6,54,0,6,44,0,3,44,2,1,162,0,2,162,3,11,163,3,1,198,0,2,306,3,2,307,3,1,337,2,3,342,0,6,334,2,6,
/* out0039_em-eta19-phi1*/	11,18,0,1,18,3,11,19,3,1,54,0,3,44,0,1,162,0,6,306,0,4,306,3,9,342,0,1,334,0,2,334,2,1,
/* out0040_em-eta0-phi2*/	0,
/* out0041_em-eta1-phi2*/	0,
/* out0042_em-eta2-phi2*/	0,
/* out0043_em-eta3-phi2*/	0,
/* out0044_em-eta4-phi2*/	3,268,1,2,272,0,5,272,1,4,
/* out0045_em-eta5-phi2*/	5,242,1,5,244,0,3,272,0,11,272,1,5,272,2,15,
/* out0046_em-eta6-phi2*/	5,208,0,1,208,1,2,242,1,5,244,0,11,244,2,8,
/* out0047_em-eta7-phi2*/	4,208,1,13,208,2,1,212,0,5,244,2,2,
/* out0048_em-eta8-phi2*/	5,176,0,5,176,1,7,208,2,2,212,0,1,212,2,3,
/* out0049_em-eta9-phi2*/	3,176,1,7,176,2,7,264,4,5,
/* out0050_em-eta10-phi2*/	9,120,4,2,142,0,9,142,1,3,264,4,11,264,5,9,265,0,14,265,1,4,265,4,1,265,5,1,
/* out0051_em-eta11-phi2*/	12,120,4,14,120,5,9,121,0,11,121,1,4,142,0,1,142,1,1,142,2,9,264,2,2,265,2,5,265,3,6,265,4,15,265,5,4,
/* out0052_em-eta12-phi2*/	13,106,1,1,110,0,6,142,2,2,120,2,2,121,0,3,121,2,4,121,3,4,121,4,16,121,5,5,234,4,6,235,1,13,265,2,4,265,3,6,
/* out0053_em-eta13-phi2*/	11,90,4,6,91,1,10,121,2,5,121,3,7,110,0,4,110,2,3,234,1,2,234,2,10,235,0,10,235,1,1,235,4,1,
/* out0054_em-eta14-phi2*/	11,74,1,2,110,2,4,90,1,2,90,2,8,91,0,10,91,1,3,91,4,1,234,2,5,234,3,6,235,3,4,235,4,5,
/* out0055_em-eta15-phi2*/	12,74,1,3,76,0,2,90,2,7,90,3,5,91,3,3,91,4,5,193,5,1,198,1,1,199,1,5,234,3,3,235,3,6,352,1,6,
/* out0056_em-eta16-phi2*/	17,44,2,1,74,1,1,76,0,2,48,5,1,49,5,1,54,1,1,55,1,4,90,3,4,91,3,8,198,1,11,198,2,1,199,1,2,337,5,1,342,1,3,343,1,6,352,1,1,352,2,6,
/* out0057_em-eta17-phi2*/	17,44,0,3,44,2,1,76,2,1,54,1,10,54,2,1,55,1,3,198,0,4,198,1,3,198,2,3,198,3,1,334,0,1,334,2,2,352,2,3,356,0,1,342,1,11,342,2,2,343,1,1,
/* out0058_em-eta18-phi2*/	13,44,0,4,54,0,4,54,1,4,54,2,3,54,3,1,198,0,3,198,3,6,334,0,5,334,2,2,342,0,5,342,1,1,342,2,2,342,3,3,
/* out0059_em-eta19-phi2*/	9,18,0,15,54,0,3,54,3,12,162,0,3,198,3,3,306,0,11,342,0,2,342,3,7,334,0,2,
/* out0060_em-eta0-phi3*/	0,
/* out0061_em-eta1-phi3*/	0,
/* out0062_em-eta2-phi3*/	0,
/* out0063_em-eta3-phi3*/	0,
/* out0064_em-eta4-phi3*/	2,272,1,1,274,0,2,
/* out0065_em-eta5-phi3*/	6,244,0,1,244,1,2,272,1,6,272,2,1,274,0,13,274,2,8,
/* out0066_em-eta6-phi3*/	5,244,0,1,244,1,14,244,2,4,248,0,5,274,2,2,
/* out0067_em-eta7-phi3*/	4,212,0,10,212,1,8,244,2,2,248,2,1,
/* out0068_em-eta8-phi3*/	4,176,1,1,178,0,3,212,1,2,212,2,12,
/* out0069_em-eta9-phi3*/	3,176,1,1,178,0,11,178,2,4,
/* out0070_em-eta10-phi3*/	7,142,1,6,146,0,1,178,2,5,264,5,7,265,5,4,270,1,2,271,1,4,
/* out0071_em-eta11-phi3*/	11,120,5,7,121,5,2,126,1,1,127,1,4,142,1,6,142,2,2,146,0,3,265,2,6,265,5,7,270,0,8,270,1,13,
/* out0072_em-eta12-phi3*/	13,110,0,4,110,1,4,146,2,1,121,2,5,121,5,9,126,0,5,126,1,14,127,1,1,234,4,10,234,5,5,265,2,1,270,0,8,270,3,3,
/* out0073_em-eta13-phi3*/	12,90,4,10,90,5,3,121,2,2,126,0,11,126,3,3,110,0,1,110,1,4,110,2,2,234,5,7,235,0,6,235,4,5,235,5,5,
/* out0074_em-eta14-phi3*/	10,76,0,1,110,2,5,90,5,10,91,0,6,91,4,4,91,5,4,235,2,8,235,3,4,235,4,5,235,5,3,
/* out0075_em-eta15-phi3*/	10,76,0,5,91,2,6,91,3,3,91,4,6,91,5,4,198,4,6,199,1,5,235,2,3,235,3,2,356,1,1,
/* out0076_em-eta16-phi3*/	13,54,4,6,55,1,4,91,2,5,91,3,2,76,0,3,76,2,2,198,2,2,199,0,8,199,1,4,342,4,6,343,1,8,356,0,5,356,1,1,
/* out0077_em-eta17-phi3*/	11,54,2,1,55,0,7,55,1,5,76,2,3,198,2,8,199,0,1,199,4,2,342,2,3,343,0,9,343,1,1,356,0,5,
/* out0078_em-eta18-phi3*/	14,44,0,2,76,2,1,54,2,8,55,0,2,55,4,2,198,2,2,198,3,3,199,3,2,199,4,2,334,0,4,356,0,1,342,2,8,342,3,1,343,4,3,
/* out0079_em-eta19-phi3*/	11,54,2,3,54,3,3,55,3,11,55,4,2,198,3,3,199,3,5,334,0,1,342,2,1,342,3,5,343,3,4,343,4,1,
/* out0080_em-eta0-phi4*/	0,
/* out0081_em-eta1-phi4*/	0,
/* out0082_em-eta2-phi4*/	0,
/* out0083_em-eta3-phi4*/	0,
/* out0084_em-eta4-phi4*/	5,274,0,1,274,1,1,292,0,11,292,1,5,292,2,8,
/* out0085_em-eta5-phi4*/	7,274,1,15,274,2,5,278,0,8,278,2,2,292,0,4,292,1,8,292,2,4,
/* out0086_em-eta6-phi4*/	5,248,0,11,248,1,11,248,2,3,274,2,1,278,2,1,
/* out0087_em-eta7-phi4*/	3,212,1,4,214,0,7,248,2,11,
/* out0088_em-eta8-phi4*/	6,178,0,1,178,1,3,212,1,2,212,2,1,214,0,5,214,2,6,
/* out0089_em-eta9-phi4*/	3,178,0,1,178,1,12,178,2,2,
/* out0090_em-eta10-phi4*/	8,146,0,6,146,1,1,178,1,1,178,2,5,270,4,12,270,5,1,271,0,1,271,1,10,
/* out0091_em-eta11-phi4*/	10,126,4,12,127,1,7,146,0,6,146,1,1,146,2,4,270,1,1,270,2,13,271,0,13,271,1,2,271,4,5,
/* out0092_em-eta12-phi4*/	13,110,1,2,146,2,6,126,1,1,126,2,11,126,5,1,127,0,13,127,1,4,127,4,4,234,5,1,270,2,3,270,3,12,271,3,9,271,4,3,
/* out0093_em-eta13-phi4*/	12,110,1,5,112,0,3,126,2,5,126,3,11,127,3,7,127,4,4,234,5,3,235,5,7,240,1,8,241,1,4,270,3,1,271,3,1,
/* out0094_em-eta14-phi4*/	16,76,0,1,76,1,1,110,1,1,110,2,1,112,0,1,112,2,1,90,5,3,91,5,6,96,1,6,97,1,4,126,3,2,127,3,3,235,2,5,235,5,1,240,0,9,240,1,4,
/* out0095_em-eta15-phi4*/	11,76,0,2,76,1,4,91,2,4,91,5,2,96,0,8,96,1,6,198,4,10,198,5,1,240,0,5,342,4,1,356,1,4,
/* out0096_em-eta16-phi4*/	12,54,4,9,91,2,1,96,0,6,76,1,2,76,2,2,198,5,7,199,0,6,342,4,9,342,5,5,356,0,1,356,1,6,356,2,1,
/* out0097_em-eta17-phi4*/	12,54,4,1,54,5,7,55,0,5,76,2,4,199,0,1,199,4,10,199,5,1,342,5,3,343,0,7,343,4,3,356,0,2,356,2,3,
/* out0098_em-eta18-phi4*/	13,55,0,2,55,4,9,55,5,1,76,2,1,199,2,2,199,3,5,199,4,2,343,2,1,343,3,5,343,4,9,343,5,1,356,0,1,356,2,2,
/* out0099_em-eta19-phi4*/	7,55,2,2,55,3,5,55,4,3,199,2,1,199,3,4,343,2,2,343,3,7,
/* out0100_em-eta0-phi5*/	0,
/* out0101_em-eta1-phi5*/	0,
/* out0102_em-eta2-phi5*/	0,
/* out0103_em-eta3-phi5*/	0,
/* out0104_em-eta4-phi5*/	6,292,0,1,292,1,2,292,2,3,296,0,5,296,1,1,296,2,3,
/* out0105_em-eta5-phi5*/	8,278,0,8,278,1,16,278,2,6,292,1,1,292,2,1,296,0,7,296,1,7,296,2,1,
/* out0106_em-eta6-phi5*/	4,248,1,4,250,0,15,250,2,1,278,2,7,
/* out0107_em-eta7-phi5*/	6,214,0,3,214,1,9,248,1,1,248,2,1,250,0,1,250,2,7,
/* out0108_em-eta8-phi5*/	4,182,0,2,214,0,1,214,1,7,214,2,9,
/* out0109_em-eta9-phi5*/	3,182,0,13,182,2,1,214,2,1,
/* out0110_em-eta10-phi5*/	5,146,1,5,182,0,1,182,2,7,270,4,4,270,5,9,
/* out0111_em-eta11-phi5*/	9,126,4,4,126,5,6,146,1,9,146,2,1,270,5,6,271,0,2,271,2,3,271,4,7,271,5,16,
/* out0112_em-eta12-phi5*/	12,112,0,4,146,2,4,126,5,9,127,0,3,127,2,1,127,4,6,127,5,15,240,4,6,241,1,1,271,2,13,271,3,6,271,4,1,
/* out0113_em-eta13-phi5*/	11,96,4,4,127,2,15,127,3,6,127,4,2,127,5,1,112,0,7,240,1,2,240,2,1,240,4,2,241,0,7,241,1,11,
/* out0114_em-eta14-phi5*/	12,96,1,1,96,2,1,96,4,4,97,0,6,97,1,12,112,0,1,112,2,6,240,0,1,240,1,2,240,2,14,240,3,2,241,0,1,
/* out0115_em-eta15-phi5*/	12,76,1,4,112,2,1,96,0,1,96,1,3,96,2,14,96,3,1,97,0,2,198,5,1,240,0,1,240,2,1,240,3,13,356,1,1,
/* out0116_em-eta16-phi5*/	11,54,5,1,96,0,1,96,2,1,96,3,13,76,1,4,198,5,7,199,5,6,240,3,1,342,5,4,356,1,3,356,2,3,
/* out0117_em-eta17-phi5*/	10,54,5,8,55,5,5,96,3,2,76,1,1,76,2,2,199,2,3,199,5,9,342,5,4,343,5,9,356,2,6,
/* out0118_em-eta18-phi5*/	7,55,2,2,55,5,10,60,0,1,199,2,9,343,2,5,343,5,6,356,2,1,
/* out0119_em-eta19-phi5*/	4,55,2,12,60,0,1,199,2,1,343,2,8,
/* out0120_em-eta0-phi6*/	0,
/* out0121_em-eta1-phi6*/	0,
/* out0122_em-eta2-phi6*/	0,
/* out0123_em-eta3-phi6*/	0,
/* out0124_em-eta4-phi6*/	6,296,0,3,296,1,1,296,2,5,298,0,3,298,1,2,298,2,1,
/* out0125_em-eta5-phi6*/	8,280,0,16,280,1,8,280,2,6,296,0,1,296,1,7,296,2,7,298,0,1,298,1,1,
/* out0126_em-eta6-phi6*/	4,250,1,15,250,2,1,254,0,4,280,2,7,
/* out0127_em-eta7-phi6*/	6,218,0,9,218,1,3,250,1,1,250,2,7,254,0,1,254,2,1,
/* out0128_em-eta8-phi6*/	4,182,1,2,218,0,7,218,1,1,218,2,9,
/* out0129_em-eta9-phi6*/	3,182,1,13,182,2,1,218,2,1,
/* out0130_em-eta10-phi6*/	5,148,0,5,182,1,1,182,2,7,276,4,4,277,1,9,
/* out0131_em-eta11-phi6*/	9,132,4,4,133,1,6,148,0,9,148,2,1,276,0,3,276,1,16,276,2,7,277,0,2,277,1,6,
/* out0132_em-eta12-phi6*/	12,112,1,4,148,2,4,132,0,1,132,1,15,132,2,6,133,0,3,133,1,9,240,4,6,240,5,1,276,0,13,276,2,1,276,3,6,
/* out0133_em-eta13-phi6*/	11,96,4,4,132,0,15,132,1,1,132,2,2,132,3,6,112,1,7,240,4,2,240,5,11,241,0,7,241,4,1,241,5,2,
/* out0134_em-eta14-phi6*/	12,96,4,4,96,5,12,97,0,6,97,4,1,97,5,1,112,1,1,112,2,6,241,0,1,241,2,1,241,3,2,241,4,14,241,5,2,
/* out0135_em-eta15-phi6*/	12,80,0,4,112,2,1,97,0,2,97,2,1,97,3,1,97,4,14,97,5,2,205,1,1,241,2,1,241,3,13,241,4,1,358,1,1,
/* out0136_em-eta16-phi6*/	11,61,1,1,97,2,1,97,3,13,97,4,1,80,0,4,204,1,6,205,1,7,241,3,1,349,1,4,358,0,3,358,1,3,
/* out0137_em-eta17-phi6*/	10,60,1,5,61,1,8,97,3,2,80,0,1,80,2,2,204,0,3,204,1,9,348,1,9,349,1,4,358,0,6,
/* out0138_em-eta18-phi6*/	6,60,0,2,60,1,10,204,0,9,348,0,5,348,1,6,358,0,1,
/* out0139_em-eta19-phi6*/	3,60,0,10,204,0,1,348,0,8,
/* out0140_em-eta0-phi7*/	0,
/* out0141_em-eta1-phi7*/	0,
/* out0142_em-eta2-phi7*/	0,
/* out0143_em-eta3-phi7*/	0,
/* out0144_em-eta4-phi7*/	5,284,0,1,284,1,1,298,0,8,298,1,5,298,2,11,
/* out0145_em-eta5-phi7*/	7,280,1,8,280,2,2,284,0,15,284,2,5,298,0,4,298,1,8,298,2,4,
/* out0146_em-eta6-phi7*/	5,254,0,11,254,1,11,254,2,3,280,2,1,284,2,1,
/* out0147_em-eta7-phi7*/	3,218,1,7,220,0,4,254,2,11,
/* out0148_em-eta8-phi7*/	6,184,0,3,184,1,1,218,1,5,218,2,6,220,0,2,220,2,1,
/* out0149_em-eta9-phi7*/	3,184,0,12,184,1,1,184,2,2,
/* out0150_em-eta10-phi7*/	8,148,0,1,148,1,6,184,0,1,184,2,5,276,4,12,276,5,10,277,0,1,277,1,1,
/* out0151_em-eta11-phi7*/	10,132,4,12,132,5,7,148,0,1,148,1,6,148,2,4,276,2,5,276,5,2,277,0,13,277,4,13,277,5,1,
/* out0152_em-eta12-phi7*/	13,116,0,2,148,2,6,132,2,4,132,5,4,133,0,13,133,1,1,133,4,11,133,5,1,247,1,1,276,2,3,276,3,9,277,3,12,277,4,3,
/* out0153_em-eta13-phi7*/	12,112,1,3,116,0,5,132,2,4,132,3,7,133,3,11,133,4,5,240,5,4,241,5,8,246,1,7,247,1,3,276,3,1,277,3,1,
/* out0154_em-eta14-phi7*/	16,80,0,1,80,1,1,112,1,1,112,2,1,116,0,1,116,2,1,96,5,4,97,5,7,102,1,6,103,1,3,132,3,3,133,3,2,241,2,9,241,5,4,246,0,5,246,1,1,
/* out0155_em-eta15-phi7*/	11,80,0,4,80,1,2,97,2,8,97,5,6,102,0,4,102,1,2,204,4,10,205,1,1,241,2,5,348,4,1,358,1,4,
/* out0156_em-eta16-phi7*/	12,60,4,9,97,2,6,102,0,1,80,0,2,80,2,2,205,0,6,205,1,7,348,4,9,349,1,5,358,0,1,358,1,6,358,2,1,
/* out0157_em-eta17-phi7*/	12,60,4,1,61,0,5,61,1,7,80,2,4,204,1,1,204,2,10,205,0,1,348,2,3,349,0,7,349,1,3,358,0,3,358,2,2,
/* out0158_em-eta18-phi7*/	13,60,1,1,60,2,9,61,0,2,80,2,1,204,0,2,204,2,2,204,3,5,348,0,1,348,1,1,348,2,9,348,3,5,358,0,2,358,2,1,
/* out0159_em-eta19-phi7*/	7,60,0,2,60,2,3,60,3,5,204,0,1,204,3,4,348,0,2,348,3,7,
/* out0160_em-eta0-phi8*/	0,
/* out0161_em-eta1-phi8*/	0,
/* out0162_em-eta2-phi8*/	0,
/* out0163_em-eta3-phi8*/	0,
/* out0164_em-eta4-phi8*/	2,284,1,2,286,1,1,
/* out0165_em-eta5-phi8*/	7,256,0,2,256,1,1,284,1,13,284,2,8,286,0,13,286,1,1,286,2,1,
/* out0166_em-eta6-phi8*/	5,254,1,5,256,0,14,256,1,1,256,2,4,284,2,2,
/* out0167_em-eta7-phi8*/	4,220,0,8,220,1,10,254,2,1,256,2,2,
/* out0168_em-eta8-phi8*/	4,184,1,3,188,0,1,220,0,2,220,2,12,
/* out0169_em-eta9-phi8*/	3,184,1,11,184,2,4,188,0,1,
/* out0170_em-eta10-phi8*/	7,148,1,1,152,0,6,184,2,5,276,5,4,277,5,2,282,1,4,283,1,7,
/* out0171_em-eta11-phi8*/	11,132,5,4,133,5,1,138,1,2,139,1,7,148,1,3,152,0,6,152,2,2,277,2,8,277,5,13,282,0,6,282,1,7,
/* out0172_em-eta12-phi8*/	13,116,0,4,116,1,4,148,2,1,132,5,1,133,2,5,133,5,14,138,0,5,138,1,9,246,4,10,247,1,5,277,2,8,277,3,3,282,0,1,
/* out0173_em-eta13-phi8*/	12,102,4,10,103,1,3,133,2,11,133,3,3,138,0,2,116,0,4,116,1,1,116,2,2,246,1,5,246,2,5,247,0,6,247,1,7,
/* out0174_em-eta14-phi8*/	10,80,1,1,116,2,5,102,1,4,102,2,4,103,0,6,103,1,10,246,0,8,246,1,3,246,2,5,246,3,4,
/* out0175_em-eta15-phi8*/	10,80,1,5,102,0,6,102,1,4,102,2,6,102,3,3,204,4,6,204,5,5,246,0,3,246,3,2,358,1,1,
/* out0176_em-eta16-phi8*/	13,60,4,6,60,5,4,102,0,5,102,3,2,80,1,3,80,2,2,204,5,4,205,0,8,205,4,2,348,4,6,348,5,8,358,1,1,358,2,5,
/* out0177_em-eta17-phi8*/	11,60,5,5,61,0,7,61,4,1,80,2,3,204,2,2,205,0,1,205,4,8,348,5,1,349,0,9,349,4,3,358,2,5,
/* out0178_em-eta18-phi8*/	14,46,1,2,80,2,1,60,2,2,61,0,2,61,4,8,204,2,2,204,3,2,205,3,3,205,4,2,338,1,4,358,2,1,348,2,3,349,3,1,349,4,8,
/* out0179_em-eta19-phi8*/	11,60,2,2,60,3,11,61,3,3,61,4,3,204,3,5,205,3,3,338,1,1,348,2,1,348,3,4,349,3,5,349,4,1,
/* out0180_em-eta0-phi9*/	0,
/* out0181_em-eta1-phi9*/	0,
/* out0182_em-eta2-phi9*/	0,
/* out0183_em-eta3-phi9*/	0,
/* out0184_em-eta4-phi9*/	2,286,1,6,290,0,2,
/* out0185_em-eta5-phi9*/	5,256,1,3,260,0,5,286,0,3,286,1,8,286,2,15,
/* out0186_em-eta6-phi9*/	5,224,0,2,224,1,1,256,1,11,256,2,8,260,0,5,
/* out0187_em-eta7-phi9*/	4,220,1,5,224,0,13,224,2,1,256,2,2,
/* out0188_em-eta8-phi9*/	5,188,0,7,188,1,5,220,1,1,220,2,3,224,2,2,
/* out0189_em-eta9-phi9*/	3,188,0,7,188,2,7,282,4,5,
/* out0190_em-eta10-phi9*/	9,138,4,2,152,0,3,152,1,9,282,1,1,282,2,1,282,4,11,282,5,4,283,0,14,283,1,9,
/* out0191_em-eta11-phi9*/	12,138,4,14,138,5,4,139,0,11,139,1,9,152,0,1,152,1,1,152,2,9,282,0,5,282,1,4,282,2,15,282,3,6,283,4,2,
/* out0192_em-eta12-phi9*/	13,116,1,6,118,0,1,152,2,2,138,0,4,138,1,5,138,2,16,138,3,4,139,0,3,139,4,2,246,4,6,246,5,13,282,0,4,282,3,6,
/* out0193_em-eta13-phi9*/	11,102,4,6,102,5,10,138,0,5,138,3,7,116,1,4,116,2,3,246,2,1,246,5,1,247,0,10,247,4,10,247,5,2,
/* out0194_em-eta14-phi9*/	11,82,0,2,116,2,4,102,2,1,102,5,3,103,0,10,103,4,8,103,5,2,246,2,5,246,3,4,247,3,6,247,4,5,
/* out0195_em-eta15-phi9*/	11,80,1,2,82,0,3,102,2,5,102,3,3,103,3,5,103,4,7,204,5,5,205,5,1,210,1,1,246,3,6,247,3,3,
/* out0196_em-eta16-phi9*/	14,60,5,4,61,5,1,66,1,1,67,1,1,102,3,8,103,3,4,80,1,2,82,0,1,204,5,2,205,4,1,205,5,11,348,5,6,349,5,3,354,1,1,
/* out0197_em-eta17-phi9*/	15,46,1,3,80,2,1,60,5,3,61,4,1,61,5,10,205,2,4,205,3,1,205,4,3,205,5,3,338,1,1,338,2,2,358,2,1,348,5,1,349,4,2,349,5,11,
/* out0198_em-eta18-phi9*/	13,46,1,4,61,2,4,61,3,1,61,4,3,61,5,4,205,2,3,205,3,6,338,1,5,338,2,2,349,2,5,349,3,3,349,4,2,349,5,1,
/* out0199_em-eta19-phi9*/	9,24,4,15,61,2,3,61,3,12,168,4,3,205,3,3,312,4,11,349,2,2,349,3,7,338,1,2,
/* out0200_em-eta0-phi10*/	0,
/* out0201_em-eta1-phi10*/	0,
/* out0202_em-eta2-phi10*/	0,
/* out0203_em-eta3-phi10*/	0,
/* out0204_em-eta4-phi10*/	2,290,0,10,290,2,1,
/* out0205_em-eta5-phi10*/	5,260,0,4,260,1,14,262,0,1,290,0,4,290,2,13,
/* out0206_em-eta6-phi10*/	5,224,1,5,226,0,3,260,0,2,260,1,1,260,2,15,
/* out0207_em-eta7-phi10*/	5,190,0,1,224,0,1,224,1,10,224,2,9,226,0,1,
/* out0208_em-eta8-phi10*/	3,188,1,8,190,0,7,224,2,4,
/* out0209_em-eta9-phi10*/	5,154,0,4,188,1,3,188,2,8,190,0,1,282,5,1,
/* out0210_em-eta10-phi10*/	8,152,1,4,154,0,8,188,2,1,282,5,11,283,0,2,283,2,3,283,4,5,283,5,15,
/* out0211_em-eta11-phi10*/	17,118,0,3,118,1,1,152,1,2,152,2,3,154,2,1,138,5,12,139,0,2,139,2,2,139,4,3,139,5,14,252,4,1,253,1,1,282,3,1,283,2,9,283,3,12,283,4,9,283,5,1,
/* out0212_em-eta12-phi10*/	13,108,4,1,138,3,1,139,2,10,139,3,10,139,4,11,139,5,2,118,0,9,246,5,2,247,5,4,252,1,7,253,1,7,282,3,3,283,3,4,
/* out0213_em-eta13-phi10*/	16,82,1,1,116,1,1,116,2,1,118,0,2,118,2,2,102,5,3,103,5,3,108,1,6,109,1,8,138,3,4,139,3,6,247,2,8,247,4,1,247,5,10,252,0,2,252,1,2,
/* out0214_em-eta14-phi10*/	10,82,0,4,82,1,2,103,2,6,103,5,11,108,0,2,108,1,4,210,4,4,211,1,1,247,2,8,247,3,6,
/* out0215_em-eta15-phi10*/	11,66,4,4,103,2,10,103,3,5,103,4,1,82,0,5,82,2,1,210,1,4,211,1,11,247,3,1,354,4,4,355,1,5,
/* out0216_em-eta16-phi10*/	11,66,1,2,67,1,12,103,3,2,82,0,1,82,2,3,205,2,1,205,5,1,210,0,2,210,1,9,354,1,7,355,1,8,
/* out0217_em-eta17-phi10*/	13,46,1,1,46,2,4,61,5,1,66,0,1,66,1,11,169,5,1,205,2,6,210,0,5,338,2,1,349,2,2,349,5,1,354,0,4,354,1,6,
/* out0218_em-eta18-phi10*/	13,24,5,1,61,2,6,66,0,6,46,1,3,46,2,1,168,4,2,168,5,11,205,2,2,312,5,2,313,5,1,349,2,6,354,0,3,338,2,6,
/* out0219_em-eta19-phi10*/	10,24,4,1,24,5,11,25,5,1,61,2,3,168,4,6,312,4,4,312,5,9,349,2,1,338,1,2,338,2,1,
/* out0220_em-eta0-phi11*/	0,
/* out0221_em-eta1-phi11*/	0,
/* out0222_em-eta2-phi11*/	0,
/* out0223_em-eta3-phi11*/	0,
/* out0224_em-eta4-phi11*/	3,262,0,1,262,1,3,290,2,1,
/* out0225_em-eta5-phi11*/	4,262,0,14,262,1,9,262,2,9,290,2,1,
/* out0226_em-eta6-phi11*/	6,226,0,9,226,1,12,226,2,2,260,1,1,260,2,1,262,2,3,
/* out0227_em-eta7-phi11*/	4,190,0,1,190,1,7,226,0,3,226,2,10,
/* out0228_em-eta8-phi11*/	3,190,0,6,190,1,5,190,2,7,
/* out0229_em-eta9-phi11*/	3,154,0,1,154,1,9,190,2,5,
/* out0230_em-eta10-phi11*/	4,154,0,3,154,1,3,154,2,7,283,2,1,
/* out0231_em-eta11-phi11*/	7,118,1,7,154,2,4,252,4,15,252,5,4,253,0,1,253,1,2,283,2,3,
/* out0232_em-eta12-phi11*/	10,108,4,15,108,5,4,139,2,4,118,0,1,118,1,4,118,2,4,252,1,3,252,2,8,253,0,11,253,1,6,
/* out0233_em-eta13-phi11*/	10,82,1,1,118,2,6,108,1,2,108,2,6,109,0,12,109,1,8,252,0,12,252,1,4,252,2,4,252,3,4,
/* out0234_em-eta14-phi11*/	11,82,1,6,108,0,10,108,1,4,108,2,6,108,3,4,210,4,12,210,5,4,211,0,1,211,1,1,252,0,2,354,4,3,
/* out0235_em-eta15-phi11*/	12,66,4,12,66,5,4,108,0,4,82,1,2,82,2,3,210,2,3,211,0,11,211,1,3,354,4,9,354,5,4,355,0,3,355,1,2,
/* out0236_em-eta16-phi11*/	12,66,2,1,67,0,12,67,1,3,82,2,4,210,0,1,210,1,2,210,2,9,210,3,1,340,1,1,354,2,6,355,0,9,355,1,1,
/* out0237_em-eta17-phi11*/	14,46,2,4,82,2,1,66,0,1,66,1,2,66,2,11,169,5,2,210,0,8,210,3,3,340,0,1,340,1,3,354,0,3,354,1,2,354,2,6,354,3,3,
/* out0238_em-eta18-phi11*/	13,46,1,1,46,2,3,66,0,8,66,3,4,168,5,4,169,0,6,169,4,4,169,5,9,313,5,6,354,0,6,354,3,1,338,2,2,340,0,3,
/* out0239_em-eta19-phi11*/	17,24,5,4,25,0,16,25,4,12,25,5,11,46,1,1,168,4,5,168,5,1,169,0,6,169,1,2,312,4,1,312,5,5,313,0,15,313,1,16,313,4,4,313,5,5,338,1,1,338,2,2,
/* out0240_em-eta0-phi12*/	0,
/* out0241_em-eta1-phi12*/	0,
/* out0242_em-eta2-phi12*/	0,
/* out0243_em-eta3-phi12*/	0,
/* out0244_em-eta4-phi12*/	1,266,0,7,
/* out0245_em-eta5-phi12*/	6,230,0,5,230,1,7,262,1,4,262,2,4,266,0,8,266,2,8,
/* out0246_em-eta6-phi12*/	6,194,1,2,226,1,4,226,2,1,230,0,11,230,1,1,230,2,7,
/* out0247_em-eta7-phi12*/	5,190,1,1,194,0,14,194,1,4,194,2,1,226,2,3,
/* out0248_em-eta8-phi12*/	6,158,0,4,158,1,3,190,1,3,190,2,4,194,0,2,194,2,3,
/* out0249_em-eta9-phi12*/	3,154,1,2,158,0,11,158,2,1,
/* out0250_em-eta10-phi12*/	7,122,0,4,122,1,1,154,1,2,154,2,4,158,0,1,158,2,1,259,1,1,
/* out0251_em-eta11-phi12*/	7,118,1,1,122,0,9,252,5,12,253,0,1,253,5,10,258,1,2,259,1,2,
/* out0252_em-eta12-phi12*/	15,86,0,1,118,1,3,118,2,2,122,0,1,122,2,1,108,5,12,109,5,7,114,1,2,115,1,2,252,2,1,253,0,3,253,2,2,253,3,3,253,4,15,253,5,5,
/* out0253_em-eta13-phi12*/	12,86,0,6,118,2,2,108,2,1,109,0,4,109,2,1,109,3,2,109,4,14,109,5,7,252,2,3,252,3,10,253,3,9,253,4,1,
/* out0254_em-eta14-phi12*/	11,82,1,2,86,0,4,108,2,3,108,3,8,109,3,10,109,4,2,210,5,12,211,0,1,211,5,5,252,3,2,354,5,3,
/* out0255_em-eta15-phi12*/	13,50,0,1,82,1,2,82,2,2,66,5,12,67,5,4,108,3,4,211,0,3,211,4,10,211,5,2,354,5,9,355,0,2,355,4,1,355,5,6,
/* out0256_em-eta16-phi12*/	14,50,0,3,82,2,2,67,0,4,67,4,9,67,5,3,210,2,4,210,3,1,211,3,3,211,4,6,340,1,4,354,2,1,355,0,2,355,4,12,355,5,1,
/* out0257_em-eta17-phi12*/	14,46,2,1,50,0,3,66,2,4,67,3,3,67,4,7,169,2,1,210,3,10,211,3,1,340,0,1,340,1,5,354,2,3,354,3,4,355,3,3,355,4,3,
/* out0258_em-eta18-phi12*/	11,46,2,3,66,3,11,67,3,1,169,2,7,169,3,1,169,4,6,169,5,4,313,2,5,313,5,1,354,3,7,340,0,5,
/* out0259_em-eta19-phi12*/	16,25,2,8,25,3,1,25,4,4,25,5,4,46,1,1,168,1,4,168,3,4,169,0,4,169,1,8,169,4,5,313,0,1,313,2,3,313,3,5,313,4,11,313,5,3,340,0,2,
/* out0260_em-eta0-phi13*/	0,
/* out0261_em-eta1-phi13*/	0,
/* out0262_em-eta2-phi13*/	0,
/* out0263_em-eta3-phi13*/	0,
/* out0264_em-eta4-phi13*/	4,232,0,1,232,1,4,266,0,1,266,2,3,
/* out0265_em-eta5-phi13*/	5,230,1,7,232,0,15,232,1,3,232,2,4,266,2,5,
/* out0266_em-eta6-phi13*/	5,194,1,2,196,0,12,196,1,2,230,1,1,230,2,9,
/* out0267_em-eta7-phi13*/	4,160,0,3,194,1,8,194,2,8,196,0,3,
/* out0268_em-eta8-phi13*/	3,158,1,9,160,0,5,194,2,4,
/* out0269_em-eta9-phi13*/	3,158,1,4,158,2,11,258,4,1,
/* out0270_em-eta10-phi13*/	7,122,1,10,124,0,1,158,2,2,258,4,15,258,5,3,259,0,7,259,1,10,
/* out0271_em-eta11-phi13*/	13,114,4,16,114,5,4,115,0,5,115,1,8,122,0,2,122,1,2,122,2,6,253,5,1,258,0,5,258,1,14,258,2,7,259,0,2,259,1,3,
/* out0272_em-eta12-phi13*/	11,86,1,5,122,2,4,109,5,1,114,0,2,114,1,14,114,2,7,115,0,4,115,1,6,216,4,7,253,2,13,258,0,7,
/* out0273_em-eta13-phi13*/	12,72,4,5,109,2,13,109,5,1,114,0,10,86,0,3,86,1,4,86,2,1,216,4,3,217,0,1,217,1,15,253,2,1,253,3,4,
/* out0274_em-eta14-phi13*/	9,72,4,5,73,1,13,109,2,2,109,3,4,86,0,2,86,2,4,211,5,5,216,0,2,216,1,13,
/* out0275_em-eta15-phi13*/	13,50,0,1,50,1,3,86,2,1,67,5,4,72,0,1,72,1,13,73,1,2,211,2,11,211,5,4,216,0,1,344,1,1,355,2,2,355,5,7,
/* out0276_em-eta16-phi13*/	15,50,0,3,50,1,1,67,2,10,67,5,5,72,0,2,174,4,1,175,1,1,211,2,4,211,3,8,340,1,2,340,2,2,344,0,1,355,2,11,355,3,2,355,5,2,
/* out0277_em-eta17-phi13*/	15,30,4,1,67,2,5,67,3,7,50,0,3,169,2,1,174,1,1,175,1,5,210,3,1,211,3,4,318,4,1,319,1,2,355,2,2,355,3,9,340,1,1,340,2,5,
/* out0278_em-eta18-phi13*/	15,31,1,5,66,3,1,67,3,5,50,0,2,50,2,1,169,2,7,169,3,5,174,1,2,313,2,3,318,1,3,319,1,4,354,3,1,355,3,2,340,0,2,340,2,3,
/* out0279_em-eta19-phi13*/	13,25,2,8,25,3,14,30,1,3,168,1,10,168,3,10,169,1,5,169,3,6,169,4,1,313,2,5,313,3,9,313,4,1,318,1,1,340,0,2,
/* out0280_em-eta0-phi14*/	0,
/* out0281_em-eta1-phi14*/	0,
/* out0282_em-eta2-phi14*/	0,
/* out0283_em-eta3-phi14*/	0,
/* out0284_em-eta4-phi14*/	4,232,1,4,236,0,12,236,1,6,236,2,7,
/* out0285_em-eta5-phi14*/	8,196,1,1,200,0,10,200,1,2,232,1,5,232,2,12,236,0,2,236,1,7,236,2,5,
/* out0286_em-eta6-phi14*/	5,164,0,1,196,0,1,196,1,13,196,2,9,200,0,3,
/* out0287_em-eta7-phi14*/	4,160,0,1,160,1,12,164,0,2,196,2,7,
/* out0288_em-eta8-phi14*/	3,160,0,7,160,1,1,160,2,10,
/* out0289_em-eta9-phi14*/	6,124,0,7,124,1,7,158,2,1,160,2,1,258,5,4,259,5,1,
/* out0290_em-eta10-phi14*/	10,114,5,1,115,5,1,122,1,2,124,0,8,124,2,3,258,5,9,259,0,6,259,2,1,259,4,8,259,5,15,
/* out0291_em-eta11-phi14*/	14,88,0,4,88,1,1,122,1,1,122,2,4,114,5,11,115,0,6,115,2,1,115,4,6,115,5,15,258,2,9,258,3,9,259,0,1,259,3,7,259,4,8,
/* out0292_em-eta12-phi14*/	12,86,1,3,88,0,5,122,2,1,114,2,9,114,3,6,115,0,1,115,3,7,115,4,10,216,4,5,216,5,13,258,0,4,258,3,6,
/* out0293_em-eta13-phi14*/	12,72,4,5,72,5,11,114,0,4,114,3,9,86,1,4,86,2,3,216,2,3,216,4,1,216,5,1,217,0,15,217,1,1,217,4,3,
/* out0294_em-eta14-phi14*/	12,72,2,1,72,4,1,72,5,3,73,0,16,73,1,1,73,4,2,86,2,6,216,0,4,216,1,3,216,2,10,216,3,3,344,1,2,
/* out0295_em-eta15-phi14*/	10,50,1,4,86,2,1,72,0,2,72,1,3,72,2,12,72,3,2,174,4,6,211,2,1,216,0,9,344,1,8,
/* out0296_em-eta16-phi14*/	13,30,4,5,67,2,1,72,0,11,72,3,1,50,1,4,50,2,1,174,4,8,175,0,1,175,1,5,318,4,10,355,2,1,344,0,6,344,1,1,
/* out0297_em-eta17-phi14*/	14,30,4,9,31,0,1,31,1,4,50,2,3,174,1,3,174,2,1,175,0,2,175,1,5,318,4,4,319,0,2,319,1,7,322,1,1,340,2,4,344,0,1,
/* out0298_em-eta18-phi14*/	13,30,1,2,30,2,1,31,0,2,31,1,7,50,2,3,174,0,1,174,1,8,318,1,5,318,2,1,319,0,1,319,1,3,322,1,2,340,2,2,
/* out0299_em-eta19-phi14*/	12,25,3,1,30,0,14,30,1,9,168,1,2,168,3,2,169,1,1,169,3,4,174,0,3,313,3,2,318,0,3,318,1,5,322,1,2,
/* out0300_em-eta0-phi15*/	0,
/* out0301_em-eta1-phi15*/	0,
/* out0302_em-eta2-phi15*/	0,
/* out0303_em-eta3-phi15*/	0,
/* out0304_em-eta4-phi15*/	3,202,1,9,236,0,2,236,2,2,
/* out0305_em-eta5-phi15*/	9,166,0,1,200,0,2,200,1,14,200,2,9,202,0,16,202,1,1,202,2,1,236,1,3,236,2,2,
/* out0306_em-eta6-phi15*/	5,164,0,4,164,1,13,166,0,1,200,0,1,200,2,7,
/* out0307_em-eta7-phi15*/	4,128,1,2,160,1,3,164,0,9,164,2,8,
/* out0308_em-eta8-phi15*/	3,128,0,10,128,1,2,160,2,5,
/* out0309_em-eta9-phi15*/	3,124,1,9,124,2,3,128,0,3,
/* out0310_em-eta10-phi15*/	5,88,1,2,92,0,1,124,2,10,222,4,6,259,2,11,
/* out0311_em-eta11-phi15*/	8,78,4,5,115,2,9,88,0,2,88,1,9,222,4,6,223,1,14,259,2,4,259,3,9,
/* out0312_em-eta12-phi15*/	13,78,4,8,79,1,12,115,2,6,115,3,8,88,0,4,88,2,5,216,5,2,217,2,1,217,5,12,222,0,1,222,1,10,223,1,1,258,3,1,
/* out0313_em-eta13-phi15*/	17,52,0,2,52,1,3,88,0,1,88,2,2,72,5,2,73,2,1,73,5,10,78,0,1,78,1,10,79,1,3,114,3,1,115,3,1,217,2,5,217,3,3,217,4,11,217,5,4,346,1,2,
/* out0314_em-eta14-phi15*/	13,52,0,6,73,2,5,73,3,2,73,4,10,73,5,6,216,2,3,216,3,8,217,3,7,217,4,2,344,1,2,344,2,2,346,0,1,346,1,2,
/* out0315_em-eta15-phi15*/	11,50,1,1,52,0,4,72,2,3,72,3,6,73,3,8,73,4,4,174,4,1,174,5,10,216,3,5,344,1,2,344,2,5,
/* out0316_em-eta16-phi15*/	11,30,4,1,30,5,8,72,3,7,50,1,3,50,2,2,174,5,4,175,0,9,318,4,1,318,5,13,344,0,5,344,2,2,
/* out0317_em-eta17-phi15*/	11,30,5,6,31,0,8,50,2,4,174,2,7,175,0,4,175,4,1,318,5,1,319,0,11,319,4,1,322,2,4,344,0,2,
/* out0318_em-eta18-phi15*/	12,30,2,6,31,0,5,31,4,1,50,2,2,174,0,3,174,1,2,174,2,4,174,3,1,318,2,9,319,0,2,322,1,3,322,2,1,
/* out0319_em-eta19-phi15*/	10,30,0,2,30,1,2,30,2,5,30,3,5,174,0,7,318,0,5,318,1,2,318,2,2,318,3,1,322,1,3,
/* out0320_em-eta0-phi16*/	0,
/* out0321_em-eta1-phi16*/	0,
/* out0322_em-eta2-phi16*/	0,
/* out0323_em-eta3-phi16*/	0,
/* out0324_em-eta4-phi16*/	3,170,1,2,202,1,6,202,2,2,
/* out0325_em-eta5-phi16*/	6,166,0,5,166,1,14,166,2,2,170,0,5,170,1,4,202,2,13,
/* out0326_em-eta6-phi16*/	6,130,0,1,130,1,4,164,1,3,164,2,2,166,0,9,166,2,8,
/* out0327_em-eta7-phi16*/	3,128,1,4,130,0,11,164,2,6,
/* out0328_em-eta8-phi16*/	3,128,0,2,128,1,8,128,2,9,
/* out0329_em-eta9-phi16*/	4,92,0,2,92,1,7,128,0,1,128,2,6,
/* out0330_em-eta10-phi16*/	6,92,0,11,92,1,1,92,2,1,222,4,3,222,5,15,223,5,5,
/* out0331_em-eta11-phi16*/	14,56,0,1,88,1,4,88,2,3,92,0,2,92,2,1,78,4,2,78,5,13,79,5,5,222,2,8,222,4,1,222,5,1,223,0,16,223,1,1,223,4,7,
/* out0332_em-eta12-phi16*/	15,56,0,2,88,2,6,78,2,4,78,4,1,78,5,3,79,0,16,79,1,1,79,4,7,79,5,1,217,2,1,222,0,12,222,1,6,222,2,7,222,3,3,346,1,1,
/* out0333_em-eta13-phi16*/	12,52,1,7,78,0,10,78,1,6,78,2,10,78,3,3,180,4,11,181,1,1,217,2,9,222,0,2,324,4,2,346,1,10,346,2,1,
/* out0334_em-eta14-phi16*/	13,36,4,10,73,2,9,78,0,4,52,0,2,52,1,2,52,2,2,180,1,2,181,1,12,217,3,6,324,4,9,325,1,4,346,0,8,346,1,1,
/* out0335_em-eta15-phi16*/	16,36,1,1,36,4,1,37,1,12,73,2,1,73,3,6,52,0,2,52,2,3,174,5,2,175,5,9,180,1,5,319,5,1,324,1,4,325,1,9,326,1,2,344,2,4,346,0,2,
/* out0336_em-eta16-phi16*/	15,22,1,1,22,2,1,52,2,1,30,5,2,31,5,8,36,1,6,37,1,1,175,4,7,175,5,7,318,5,2,319,5,12,324,1,2,326,1,3,344,0,1,344,2,3,
/* out0337_em-eta17-phi16*/	10,22,1,3,31,4,6,31,5,8,174,2,2,175,3,1,175,4,8,319,4,10,319,5,3,322,2,5,326,0,1,
/* out0338_em-eta18-phi16*/	14,22,1,2,30,2,1,31,3,1,31,4,9,174,2,2,174,3,7,175,3,1,318,2,4,318,3,1,319,3,1,319,4,5,322,0,2,322,1,1,322,2,3,
/* out0339_em-eta19-phi16*/	8,30,2,3,30,3,7,31,3,1,174,0,2,174,3,3,318,0,8,318,3,9,322,1,3,
/* out0340_em-eta0-phi17*/	0,
/* out0341_em-eta1-phi17*/	0,
/* out0342_em-eta2-phi17*/	0,
/* out0343_em-eta3-phi17*/	0,
/* out0344_em-eta4-phi17*/	1,170,1,4,
/* out0345_em-eta5-phi17*/	7,134,0,4,134,1,8,166,1,2,166,2,3,170,0,11,170,1,6,170,2,16,
/* out0346_em-eta6-phi17*/	4,130,1,10,130,2,1,134,0,12,166,2,3,
/* out0347_em-eta7-phi17*/	4,94,1,1,130,0,3,130,1,2,130,2,15,
/* out0348_em-eta8-phi17*/	4,94,0,9,94,1,7,128,2,1,130,0,1,
/* out0349_em-eta9-phi17*/	3,92,1,7,92,2,1,94,0,7,
/* out0350_em-eta10-phi17*/	4,92,1,1,92,2,11,223,2,5,223,5,8,
/* out0351_em-eta11-phi17*/	11,56,0,1,56,1,7,92,2,2,79,2,3,79,5,6,223,2,11,223,3,11,223,4,9,223,5,3,350,0,3,350,1,3,
/* out0352_em-eta12-phi17*/	16,56,0,8,56,1,1,79,2,13,79,3,8,79,4,8,79,5,4,180,4,1,180,5,6,222,0,1,222,2,1,222,3,13,223,3,5,346,2,1,350,0,13,350,1,1,350,2,7,
/* out0353_em-eta13-phi17*/	16,36,5,4,78,0,1,78,2,2,78,3,13,79,3,8,79,4,1,52,1,4,56,0,4,180,4,4,180,5,10,181,0,9,181,1,1,324,4,2,324,5,11,346,2,10,350,2,1,
/* out0354_em-eta14-phi17*/	15,36,4,5,36,5,12,37,0,7,52,2,6,180,1,2,180,2,7,181,0,7,181,1,2,324,4,3,324,5,5,325,0,13,325,1,2,326,1,1,346,0,5,346,2,4,
/* out0355_em-eta15-phi17*/	15,22,2,1,52,2,4,36,1,1,36,2,7,37,0,9,37,1,3,175,2,1,180,0,7,180,1,7,180,2,1,324,1,6,324,2,8,325,0,3,325,1,1,326,1,7,
/* out0356_em-eta16-phi17*/	11,22,2,5,36,0,6,36,1,8,36,2,1,175,2,13,180,0,1,319,2,4,324,0,8,324,1,4,326,0,3,326,1,3,
/* out0357_em-eta17-phi17*/	9,22,1,3,31,2,12,36,0,2,175,2,2,175,3,9,319,2,12,319,3,2,322,2,2,326,0,4,
/* out0358_em-eta18-phi17*/	8,22,1,2,31,2,4,31,3,8,174,3,4,175,3,5,319,3,10,322,0,8,322,2,1,
/* out0359_em-eta19-phi17*/	7,30,3,4,31,3,6,174,3,1,318,3,5,319,3,3,322,0,6,322,1,1,
/* out0360_em-eta0-phi18*/	0,
/* out0361_em-eta1-phi18*/	0,
/* out0362_em-eta2-phi18*/	0,
/* out0363_em-eta3-phi18*/	0,
/* out0364_em-eta4-phi18*/	1,136,1,5,
/* out0365_em-eta5-phi18*/	7,100,0,3,100,1,2,134,1,8,134,2,4,136,0,16,136,1,10,136,2,9,
/* out0366_em-eta6-phi18*/	4,98,0,1,98,1,10,100,0,3,134,2,12,
/* out0367_em-eta7-phi18*/	4,94,1,1,98,0,15,98,1,2,98,2,3,
/* out0368_em-eta8-phi18*/	4,62,0,1,94,1,7,94,2,9,98,2,1,
/* out0369_em-eta9-phi18*/	3,58,0,1,58,1,7,94,2,7,
/* out0370_em-eta10-phi18*/	4,58,0,11,58,1,1,186,4,5,186,5,8,
/* out0371_em-eta11-phi18*/	14,42,4,3,42,5,6,56,1,7,56,2,1,58,0,2,186,4,11,186,5,3,187,0,9,187,1,11,330,4,11,330,5,10,331,0,1,332,0,1,350,1,5,
/* out0372_em-eta12-phi18*/	20,42,4,13,42,5,4,43,0,8,43,1,8,56,1,1,56,2,8,181,2,1,181,5,6,186,0,1,186,1,13,186,2,1,187,1,5,328,1,1,350,1,7,350,2,6,330,1,2,330,2,2,330,4,5,331,0,8,331,1,15,
/* out0373_em-eta13-phi18*/	19,26,1,4,56,2,4,37,5,4,42,0,1,42,1,13,42,2,2,43,0,1,43,1,8,181,2,4,181,3,1,181,4,9,181,5,10,325,2,2,325,5,11,330,0,1,330,1,11,331,1,1,328,1,10,350,2,2,
/* out0374_em-eta14-phi18*/	15,26,0,6,37,2,5,37,4,7,37,5,12,180,2,7,180,3,2,181,3,2,181,4,7,325,2,3,325,3,2,325,4,13,325,5,5,326,2,1,328,0,5,328,1,4,
/* out0375_em-eta15-phi18*/	15,22,2,1,26,0,4,36,2,7,36,3,1,37,3,3,37,4,9,144,4,1,180,0,7,180,2,1,180,3,7,324,2,8,324,3,6,325,3,1,325,4,3,326,2,7,
/* out0376_em-eta16-phi18*/	11,22,2,5,36,0,6,36,2,1,36,3,8,144,4,13,180,0,1,288,4,4,324,0,8,324,3,4,326,0,3,326,2,3,
/* out0377_em-eta17-phi18*/	11,0,4,12,36,0,2,22,0,3,22,1,2,22,2,1,144,4,2,145,1,9,288,4,12,289,1,2,310,2,2,326,0,4,
/* out0378_em-eta18-phi18*/	8,0,4,4,1,1,8,22,1,2,144,1,4,145,1,5,289,1,10,310,1,3,310,2,1,
/* out0379_em-eta19-phi18*/	6,0,1,4,1,1,6,144,1,1,288,1,5,289,1,3,310,1,3,
/* out0380_em-eta0-phi19*/	0,
/* out0381_em-eta1-phi19*/	0,
/* out0382_em-eta2-phi19*/	0,
/* out0383_em-eta3-phi19*/	0,
/* out0384_em-eta4-phi19*/	3,104,1,8,136,1,1,136,2,1,
/* out0385_em-eta5-phi19*/	7,100,0,2,100,1,14,100,2,5,104,0,16,104,1,5,104,2,2,136,2,6,
/* out0386_em-eta6-phi19*/	6,64,0,2,64,1,3,98,1,4,98,2,1,100,0,8,100,2,9,
/* out0387_em-eta7-phi19*/	3,62,1,4,64,0,6,98,2,11,
/* out0388_em-eta8-phi19*/	3,62,0,9,62,1,8,62,2,2,
/* out0389_em-eta9-phi19*/	4,58,1,7,58,2,2,62,0,6,62,2,1,
/* out0390_em-eta10-phi19*/	6,58,0,1,58,1,1,58,2,11,186,5,5,187,2,3,187,5,15,
/* out0391_em-eta11-phi19*/	21,28,0,3,28,1,4,56,2,1,58,0,1,58,2,2,42,5,5,43,2,2,43,5,13,186,2,8,187,0,7,187,2,1,187,3,1,187,4,16,187,5,1,330,5,6,331,0,2,331,2,4,331,4,5,331,5,16,332,0,3,332,1,5,
/* out0392_em-eta12-phi19*/	23,28,0,6,56,2,2,42,2,4,42,5,1,43,0,7,43,2,1,43,3,1,43,4,16,43,5,3,150,4,1,186,0,12,186,1,3,186,2,7,186,3,6,328,2,1,332,0,12,332,1,1,332,2,7,330,2,13,330,3,2,331,0,5,331,3,1,331,4,11,
/* out0393_em-eta13-phi19*/	17,26,1,7,42,0,10,42,1,3,42,2,10,42,3,6,150,4,9,181,2,11,181,3,1,186,0,2,294,4,3,325,2,2,330,0,14,330,1,3,330,2,1,330,3,4,328,1,1,328,2,10,
/* out0394_em-eta14-phi19*/	15,6,4,9,37,2,10,42,0,4,26,0,2,26,1,2,26,2,2,151,1,6,180,3,2,181,3,12,294,4,7,295,1,2,325,2,9,325,3,4,328,0,8,328,2,1,
/* out0395_em-eta15-phi19*/	17,6,4,1,7,1,6,36,3,1,37,2,1,37,3,12,26,0,3,26,2,2,144,5,9,145,5,2,180,3,5,288,5,1,295,1,4,324,3,4,325,3,9,314,1,4,326,2,2,328,0,2,
/* out0396_em-eta16-phi19*/	15,0,5,8,1,5,2,36,3,6,37,3,1,22,0,3,22,2,2,26,0,1,144,5,7,145,0,7,288,5,12,289,5,2,324,3,2,314,0,1,314,1,3,326,2,3,
/* out0397_em-eta17-phi19*/	10,0,5,8,1,0,6,22,0,8,144,2,2,145,0,8,145,1,1,288,5,3,289,0,10,310,2,5,326,0,1,
/* out0398_em-eta18-phi19*/	14,0,2,1,1,0,9,1,1,1,22,0,1,22,1,1,144,1,7,144,2,2,145,1,1,288,1,1,288,2,4,289,0,5,289,1,1,310,1,2,310,2,3,
/* out0399_em-eta19-phi19*/	8,0,1,7,0,2,3,1,1,1,144,0,2,144,1,3,288,0,8,288,1,9,310,1,3,
/* out0400_em-eta0-phi20*/	0,
/* out0401_em-eta1-phi20*/	0,
/* out0402_em-eta2-phi20*/	0,
/* out0403_em-eta3-phi20*/	0,
/* out0404_em-eta4-phi20*/	4,70,0,2,70,2,2,104,1,3,104,2,6,
/* out0405_em-eta5-phi20*/	7,68,0,9,68,1,14,68,2,2,70,0,2,70,1,3,100,2,1,104,2,8,
/* out0406_em-eta6-phi20*/	5,64,1,13,64,2,4,68,0,7,68,2,1,100,2,1,
/* out0407_em-eta7-phi20*/	4,34,1,3,62,1,2,64,0,8,64,2,9,
/* out0408_em-eta8-phi20*/	3,34,0,5,62,1,2,62,2,10,
/* out0409_em-eta9-phi20*/	3,32,0,3,32,1,9,62,2,3,
/* out0410_em-eta10-phi20*/	5,28,1,2,32,0,10,58,2,1,156,4,11,187,2,6,
/* out0411_em-eta11-phi20*/	13,12,4,9,43,2,5,28,1,9,28,2,2,156,4,4,157,1,9,187,2,6,187,3,14,300,4,14,301,1,1,331,2,11,320,0,2,332,1,7,
/* out0412_em-eta12-phi20*/	23,12,4,6,13,1,8,43,2,8,43,3,12,28,0,5,28,2,4,150,4,1,150,5,12,151,5,2,156,1,1,186,0,1,186,3,10,187,3,1,295,5,1,300,1,1,300,4,1,301,1,8,330,3,5,331,2,1,331,3,15,316,1,2,332,1,3,332,2,8,
/* out0413_em-eta13-phi20*/	25,6,4,1,6,5,10,7,5,2,12,1,1,13,1,1,42,0,1,42,3,10,43,3,3,26,1,3,26,2,2,28,0,2,28,2,1,150,4,5,150,5,4,151,0,11,151,1,3,294,4,3,294,5,15,295,0,2,295,5,2,330,0,1,330,3,5,316,1,8,328,2,2,332,2,1,
/* out0414_em-eta14-phi20*/	20,6,4,5,6,5,6,7,0,10,7,1,2,26,2,6,150,1,8,150,2,3,151,0,2,151,1,7,294,2,1,294,4,3,294,5,1,295,0,12,295,1,6,314,1,2,314,2,2,316,0,2,316,1,2,328,0,1,328,2,2,
/* out0415_em-eta15-phi20*/	14,2,1,1,26,2,4,6,1,6,6,2,3,7,0,4,7,1,8,145,2,1,145,5,10,150,1,5,294,1,12,294,2,2,295,1,4,314,1,5,314,2,2,
/* out0416_em-eta16-phi20*/	12,1,2,1,1,5,8,6,1,7,2,0,2,2,1,3,145,4,9,145,5,4,289,2,1,289,5,13,294,1,1,314,0,5,314,1,2,
/* out0417_em-eta17-phi20*/	11,1,4,8,1,5,6,2,0,4,144,2,7,145,0,1,145,4,4,289,0,1,289,4,11,289,5,1,310,2,4,314,0,2,
/* out0418_em-eta18-phi20*/	14,0,2,6,1,0,1,1,4,5,2,0,2,22,0,1,144,0,3,144,1,1,144,2,4,144,3,2,288,2,9,289,4,2,310,0,7,310,1,1,310,2,1,
/* out0419_em-eta19-phi20*/	10,0,0,2,0,1,5,0,2,5,0,3,2,144,0,7,288,0,5,288,1,1,288,2,2,288,3,2,310,1,3,
/* out0420_em-eta0-phi21*/	0,
/* out0421_em-eta1-phi21*/	0,
/* out0422_em-eta2-phi21*/	0,
/* out0423_em-eta3-phi21*/	0,
/* out0424_em-eta4-phi21*/	4,40,1,4,70,0,7,70,1,6,70,2,12,
/* out0425_em-eta5-phi21*/	8,38,1,1,40,0,12,40,1,5,68,1,2,68,2,10,70,0,5,70,1,7,70,2,2,
/* out0426_em-eta6-phi21*/	5,38,0,9,38,1,13,38,2,1,64,2,1,68,2,3,
/* out0427_em-eta7-phi21*/	4,34,1,12,34,2,1,38,0,7,64,2,2,
/* out0428_em-eta8-phi21*/	3,34,0,10,34,1,1,34,2,7,
/* out0429_em-eta9-phi21*/	6,10,0,1,32,1,7,32,2,7,34,0,1,156,5,1,157,5,4,
/* out0430_em-eta10-phi21*/	12,8,1,2,32,0,3,32,2,8,12,5,1,13,5,1,156,4,1,156,5,15,157,0,8,157,4,6,157,5,9,300,5,6,301,5,9,
/* out0431_em-eta11-phi21*/	23,8,0,4,8,1,1,28,1,1,28,2,4,12,4,1,12,5,15,13,0,6,13,4,6,13,5,11,156,1,9,156,2,9,157,0,8,157,1,7,157,4,1,300,2,2,300,4,1,300,5,10,301,0,14,301,1,2,301,4,7,301,5,3,320,0,10,320,2,1,
/* out0432_em-eta12-phi21*/	21,4,1,3,8,0,1,28,2,5,12,1,6,12,2,9,13,0,10,13,1,7,13,4,1,151,2,5,151,5,13,156,0,4,156,1,6,300,0,2,300,1,15,300,2,7,301,0,2,301,1,5,316,1,1,316,2,6,320,0,2,320,2,7,
/* out0433_em-eta13-phi21*/	19,4,0,3,4,1,4,7,2,5,7,5,11,12,0,4,12,1,9,150,2,3,151,0,3,151,2,1,151,3,1,151,4,15,151,5,1,295,2,6,295,4,5,295,5,13,300,0,1,316,0,4,316,1,3,316,2,5,
/* out0434_em-eta14-phi21*/	17,4,0,6,6,2,1,7,0,2,7,2,1,7,3,1,7,4,16,7,5,3,150,0,4,150,1,3,150,2,10,150,3,3,294,2,8,295,0,2,295,3,1,295,4,11,314,2,2,316,0,7,
/* out0435_em-eta15-phi21*/	13,2,1,4,4,0,1,6,0,2,6,1,2,6,2,12,6,3,3,145,2,6,150,0,9,294,0,8,294,1,3,294,2,5,294,3,3,314,2,8,
/* out0436_em-eta16-phi21*/	12,1,2,5,6,0,11,6,1,1,2,0,1,2,1,4,145,2,8,145,3,5,145,4,1,289,2,10,294,0,5,314,0,6,314,2,1,
/* out0437_em-eta17-phi21*/	14,1,2,9,1,3,4,1,4,1,2,0,3,144,2,1,144,3,3,145,3,5,145,4,2,289,2,4,289,3,7,289,4,2,302,1,4,310,0,1,314,0,1,
/* out0438_em-eta18-phi21*/	13,0,2,1,0,3,2,1,3,7,1,4,2,2,0,3,144,0,1,144,3,8,288,2,1,288,3,5,289,3,3,289,4,1,302,1,2,310,0,6,
/* out0439_em-eta19-phi21*/	8,0,0,14,0,3,9,144,0,3,288,0,3,288,3,5,302,0,1,310,0,2,310,1,1,
/* out0440_em-eta0-phi22*/	0,
/* out0441_em-eta1-phi22*/	0,
/* out0442_em-eta2-phi22*/	0,
/* out0443_em-eta3-phi22*/	0,
/* out0444_em-eta4-phi22*/	3,20,0,4,40,1,4,40,2,1,
/* out0445_em-eta5-phi22*/	6,16,1,7,20,0,5,20,2,1,40,0,4,40,1,3,40,2,15,
/* out0446_em-eta6-phi22*/	5,14,1,2,16,0,9,16,1,1,38,1,2,38,2,12,
/* out0447_em-eta7-phi22*/	4,14,0,8,14,1,8,34,2,3,38,2,3,
/* out0448_em-eta8-phi22*/	3,10,1,9,14,0,4,34,2,5,
/* out0449_em-eta9-phi22*/	3,10,0,11,10,1,4,157,2,1,
/* out0450_em-eta10-phi22*/	9,8,1,10,10,0,2,32,2,1,157,2,15,157,3,10,157,4,7,157,5,3,301,2,8,301,5,2,
/* out0451_em-eta11-phi22*/	22,8,0,6,8,1,2,8,2,2,13,2,16,13,3,8,13,4,5,13,5,4,156,0,5,156,2,7,156,3,14,157,3,3,157,4,2,300,2,2,300,3,1,301,2,8,301,3,13,301,4,9,301,5,2,308,1,1,308,2,3,320,0,2,320,2,3,
/* out0452_em-eta12-phi22*/	15,4,1,5,8,0,4,12,0,2,12,2,7,12,3,14,13,3,6,13,4,4,151,2,7,156,0,7,300,0,10,300,2,5,300,3,13,308,1,8,316,2,1,320,2,5,
/* out0453_em-eta13-phi22*/	16,4,0,1,4,1,4,4,2,3,7,2,5,12,0,10,151,2,3,151,3,15,151,4,1,295,2,10,295,3,1,300,0,3,304,2,1,308,0,1,308,1,4,316,0,2,316,2,4,
/* out0454_em-eta14-phi22*/	11,4,0,4,4,2,2,7,2,5,7,3,13,150,0,2,150,3,13,294,3,5,295,3,14,304,1,8,304,2,1,316,0,1,
/* out0455_em-eta15-phi22*/	12,2,1,3,2,2,1,4,0,1,6,0,1,6,3,13,7,3,2,150,0,1,294,0,3,294,3,8,304,0,2,304,1,6,314,2,1,
/* out0456_em-eta16-phi22*/	9,2,1,1,2,2,3,6,0,2,145,2,1,145,3,1,302,1,2,302,2,3,304,0,2,314,0,1,
/* out0457_em-eta17-phi22*/	9,1,2,1,2,2,3,144,3,1,145,3,5,289,2,1,289,3,2,302,0,1,302,1,5,302,2,1,
/* out0458_em-eta18-phi22*/	8,1,3,5,2,0,1,2,2,2,144,3,2,288,3,3,289,3,4,302,0,2,302,1,3,
/* out0459_em-eta19-phi22*/	3,0,3,3,288,3,1,302,0,3,
/* out0460_em-eta0-phi23*/	0,
/* out0461_em-eta1-phi23*/	0,
/* out0462_em-eta2-phi23*/	0,
/* out0463_em-eta3-phi23*/	0,
/* out0464_em-eta4-phi23*/	2,20,0,5,20,2,1,
/* out0465_em-eta5-phi23*/	4,16,1,7,16,2,5,20,0,2,20,2,14,
/* out0466_em-eta6-phi23*/	4,14,1,2,16,0,7,16,1,1,16,2,11,
/* out0467_em-eta7-phi23*/	3,14,0,1,14,1,4,14,2,14,
/* out0468_em-eta8-phi23*/	4,10,1,3,10,2,4,14,0,3,14,2,2,
/* out0469_em-eta9-phi23*/	2,10,0,1,10,2,11,
/* out0470_em-eta10-phi23*/	5,8,1,1,8,2,4,10,0,1,10,2,1,157,3,1,
/* out0471_em-eta11-phi23*/	5,8,2,9,156,3,2,157,3,2,301,3,3,308,2,4,
/* out0472_em-eta12-phi23*/	9,4,2,1,8,0,1,8,2,1,12,3,2,13,3,2,300,3,2,308,0,6,308,1,3,308,2,9,
/* out0473_em-eta13-phi23*/	3,4,2,6,304,2,2,308,0,9,
/* out0474_em-eta14-phi23*/	4,4,2,4,304,0,1,304,1,1,304,2,9,
/* out0475_em-eta15-phi23*/	4,2,2,1,304,0,8,304,1,1,304,2,3,
/* out0476_em-eta16-phi23*/	3,2,2,3,302,2,7,304,0,3,
/* out0477_em-eta17-phi23*/	3,2,2,3,302,0,1,302,2,5,
/* out0478_em-eta18-phi23*/	1,302,0,5,
/* out0479_em-eta19-phi23*/	1,302,0,3
};
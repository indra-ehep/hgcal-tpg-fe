parameter integer matrixH [0:11282] = {
/* num inputs = 360(in0-in359) */
/* num outputs = 600(out0-out599) */
//* max inputs per outputs = 25 */
//* total number of input in adders 3560 */

/* out0000_em-eta0-phi0*/	0,
/* out0001_em-eta1-phi0*/	0,
/* out0002_em-eta2-phi0*/	0,
/* out0003_em-eta3-phi0*/	0,
/* out0004_em-eta4-phi0*/	0,
/* out0005_em-eta5-phi0*/	0,
/* out0006_em-eta6-phi0*/	0,
/* out0007_em-eta7-phi0*/	0,
/* out0008_em-eta8-phi0*/	0,
/* out0009_em-eta9-phi0*/	0,
/* out0010_em-eta10-phi0*/	0,
/* out0011_em-eta11-phi0*/	0,
/* out0012_em-eta12-phi0*/	0,
/* out0013_em-eta13-phi0*/	0,
/* out0014_em-eta14-phi0*/	0,
/* out0015_em-eta15-phi0*/	0,
/* out0016_em-eta16-phi0*/	0,
/* out0017_em-eta17-phi0*/	0,
/* out0018_em-eta18-phi0*/	0,
/* out0019_em-eta19-phi0*/	0,
/* out0020_em-eta0-phi1*/	0,
/* out0021_em-eta1-phi1*/	0,
/* out0022_em-eta2-phi1*/	0,
/* out0023_em-eta3-phi1*/	0,
/* out0024_em-eta4-phi1*/	0,
/* out0025_em-eta5-phi1*/	0,
/* out0026_em-eta6-phi1*/	0,
/* out0027_em-eta7-phi1*/	0,
/* out0028_em-eta8-phi1*/	0,
/* out0029_em-eta9-phi1*/	0,
/* out0030_em-eta10-phi1*/	0,
/* out0031_em-eta11-phi1*/	0,
/* out0032_em-eta12-phi1*/	0,
/* out0033_em-eta13-phi1*/	0,
/* out0034_em-eta14-phi1*/	0,
/* out0035_em-eta15-phi1*/	1,36,0,1,
/* out0036_em-eta16-phi1*/	2,42,0,1,38,0,1,
/* out0037_em-eta17-phi1*/	0,
/* out0038_em-eta18-phi1*/	0,
/* out0039_em-eta19-phi1*/	6,19,5,1,16,1,1,16,5,2,17,1,2,17,5,4,17,5,2,
/* out0040_em-eta0-phi2*/	0,
/* out0041_em-eta1-phi2*/	0,
/* out0042_em-eta2-phi2*/	0,
/* out0043_em-eta3-phi2*/	0,
/* out0044_em-eta4-phi2*/	0,
/* out0045_em-eta5-phi2*/	0,
/* out0046_em-eta6-phi2*/	0,
/* out0047_em-eta7-phi2*/	0,
/* out0048_em-eta8-phi2*/	0,
/* out0049_em-eta9-phi2*/	0,
/* out0050_em-eta10-phi2*/	0,
/* out0051_em-eta11-phi2*/	1,60,1,1,
/* out0052_em-eta12-phi2*/	2,68,1,1,60,0,13,
/* out0053_em-eta13-phi2*/	4,68,0,13,68,1,1,60,0,1,60,3,4,
/* out0054_em-eta14-phi2*/	3,68,0,2,68,3,4,36,1,5,
/* out0055_em-eta15-phi2*/	5,42,1,4,36,0,11,36,1,4,38,0,2,38,1,7,
/* out0056_em-eta16-phi2*/	7,42,0,10,42,1,5,36,0,4,36,3,8,38,0,11,38,1,2,38,3,2,
/* out0057_em-eta17-phi2*/	7,42,0,5,42,3,7,17,2,1,36,3,4,37,3,1,38,0,2,38,3,9,
/* out0058_em-eta18-phi2*/	7,42,3,5,43,3,1,17,2,7,17,5,5,17,2,3,38,3,2,39,3,1,
/* out0059_em-eta19-phi2*/	10,19,2,8,19,5,14,16,1,5,16,5,10,17,1,10,17,4,1,17,5,6,17,2,5,17,4,1,17,5,9,
/* out0060_em-eta0-phi3*/	0,
/* out0061_em-eta1-phi3*/	0,
/* out0062_em-eta2-phi3*/	0,
/* out0063_em-eta3-phi3*/	0,
/* out0064_em-eta4-phi3*/	0,
/* out0065_em-eta5-phi3*/	2,158,0,4,158,2,4,
/* out0066_em-eta6-phi3*/	2,136,0,4,136,2,1,
/* out0067_em-eta7-phi3*/	2,114,0,1,136,2,3,
/* out0068_em-eta8-phi3*/	2,114,0,3,114,2,4,
/* out0069_em-eta9-phi3*/	1,92,0,2,
/* out0070_em-eta10-phi3*/	2,92,0,2,92,2,4,
/* out0071_em-eta11-phi3*/	4,70,0,1,60,1,10,61,0,1,61,1,12,
/* out0072_em-eta12-phi3*/	10,68,1,7,69,1,12,70,0,3,70,2,2,60,0,2,60,1,5,60,2,15,60,3,3,61,0,3,61,4,1,
/* out0073_em-eta13-phi3*/	11,68,0,1,68,1,7,68,2,14,68,3,2,69,0,4,69,4,1,70,2,2,60,2,1,60,3,9,61,3,10,61,4,3,
/* out0074_em-eta14-phi3*/	10,48,0,2,68,2,2,68,3,10,69,3,8,69,4,3,36,1,5,37,0,1,37,1,12,61,3,2,39,1,3,
/* out0075_em-eta15-phi3*/	12,42,1,4,43,1,12,69,3,4,48,0,2,48,2,2,36,1,2,36,2,10,37,0,3,38,1,6,38,2,1,39,0,2,39,1,9,
/* out0076_em-eta16-phi3*/	12,42,1,3,42,2,9,43,0,4,48,2,2,36,2,6,36,3,3,37,3,1,37,4,4,38,1,1,38,2,12,39,0,2,39,4,1,
/* out0077_em-eta17-phi3*/	11,28,2,1,42,2,7,42,3,3,43,4,4,17,2,1,36,3,1,37,3,10,38,2,3,38,3,3,39,3,4,39,4,3,
/* out0078_em-eta18-phi3*/	10,28,2,3,42,3,1,43,3,11,17,2,7,17,3,4,17,4,6,17,5,1,17,2,5,17,3,1,39,3,7,
/* out0079_em-eta19-phi3*/	15,19,2,8,19,3,4,19,4,4,19,5,1,28,0,1,16,1,8,16,2,4,16,5,4,17,1,4,17,4,5,16,2,1,17,2,3,17,3,3,17,4,11,17,5,5,
/* out0080_em-eta0-phi4*/	0,
/* out0081_em-eta1-phi4*/	0,
/* out0082_em-eta2-phi4*/	0,
/* out0083_em-eta3-phi4*/	0,
/* out0084_em-eta4-phi4*/	3,158,0,3,158,1,1,178,2,2,
/* out0085_em-eta5-phi4*/	4,158,0,9,158,1,14,158,2,9,178,2,1,
/* out0086_em-eta6-phi4*/	6,136,0,12,136,1,9,136,2,2,158,2,3,160,0,1,160,2,1,
/* out0087_em-eta7-phi4*/	4,114,0,7,114,1,1,136,1,3,136,2,10,
/* out0088_em-eta8-phi4*/	3,114,0,5,114,1,6,114,2,7,
/* out0089_em-eta9-phi4*/	3,92,0,9,92,1,1,114,2,5,
/* out0090_em-eta10-phi4*/	4,92,0,3,92,1,3,92,2,7,86,0,1,
/* out0091_em-eta11-phi4*/	7,70,0,7,92,2,4,60,4,15,60,5,2,61,0,1,61,1,4,86,0,3,
/* out0092_em-eta12-phi4*/	10,68,4,15,69,1,4,96,0,4,70,0,4,70,1,1,70,2,4,60,5,6,61,0,11,61,4,8,61,5,3,
/* out0093_em-eta13-phi4*/	10,48,0,1,70,2,6,68,5,8,69,0,12,69,4,6,69,5,2,61,2,12,61,3,4,61,4,4,61,5,4,
/* out0094_em-eta14-phi4*/	11,48,0,6,69,2,10,69,3,4,69,4,6,69,5,4,36,4,12,36,5,1,37,0,1,37,1,4,61,2,2,38,4,3,
/* out0095_em-eta15-phi4*/	13,42,4,12,43,1,4,69,2,4,48,0,2,48,2,3,36,5,3,37,0,11,37,4,3,38,4,9,38,5,2,39,0,3,39,1,4,234,0,4,
/* out0096_em-eta16-phi4*/	12,42,5,3,43,0,12,43,4,1,48,2,4,37,2,1,37,3,1,37,4,9,37,5,2,38,5,1,39,0,9,39,4,6,234,0,5,
/* out0097_em-eta17-phi4*/	13,28,2,4,48,2,1,43,2,1,43,4,11,43,5,2,17,3,2,37,2,8,37,3,3,39,2,3,39,3,3,39,4,6,39,5,2,234,0,2,
/* out0098_em-eta18-phi4*/	12,28,0,1,28,2,3,43,2,8,43,3,4,16,2,6,16,3,4,17,3,9,17,4,4,17,3,6,39,2,6,39,3,1,222,2,2,
/* out0099_em-eta19-phi4*/	17,18,2,16,18,3,4,19,3,11,19,4,12,28,0,1,16,0,5,16,1,2,16,2,6,16,3,1,16,0,1,16,1,16,16,2,15,16,3,5,17,3,5,17,4,4,222,0,1,222,2,2,
/* out0100_em-eta0-phi5*/	0,
/* out0101_em-eta1-phi5*/	0,
/* out0102_em-eta2-phi5*/	0,
/* out0103_em-eta3-phi5*/	0,
/* out0104_em-eta4-phi5*/	2,178,1,3,178,2,8,
/* out0105_em-eta5-phi5*/	5,158,1,1,160,0,14,160,1,4,178,1,11,178,2,5,
/* out0106_em-eta6-phi5*/	5,136,1,3,138,0,5,160,0,1,160,1,2,160,2,15,
/* out0107_em-eta7-phi5*/	5,114,1,1,136,1,1,138,0,10,138,1,1,138,2,9,
/* out0108_em-eta8-phi5*/	3,114,1,7,116,0,8,138,2,4,
/* out0109_em-eta9-phi5*/	5,92,1,4,114,1,1,116,0,3,116,2,8,87,1,1,
/* out0110_em-eta10-phi5*/	8,92,1,8,94,0,4,116,2,1,86,0,3,86,1,15,86,2,5,87,0,2,87,1,11,
/* out0111_em-eta11-phi5*/	17,70,0,1,70,1,3,92,2,1,94,0,2,94,2,3,96,0,2,96,1,14,96,2,3,97,0,2,97,1,12,60,4,1,60,5,1,86,0,9,86,1,1,86,2,9,86,3,12,87,3,1,
/* out0112_em-eta12-phi5*/	13,68,4,1,96,0,10,96,1,2,96,2,11,96,3,10,97,3,1,70,1,9,60,5,7,61,5,7,62,1,4,63,1,2,86,3,4,87,3,3,
/* out0113_em-eta13-phi5*/	16,48,0,1,70,1,2,70,2,2,72,0,1,72,2,1,68,5,8,69,5,6,70,1,3,71,1,3,96,3,6,97,3,4,61,2,2,61,5,2,62,0,8,62,1,10,62,2,1,
/* out0114_em-eta14-phi5*/	11,48,0,2,48,1,4,69,2,2,69,5,4,70,0,6,70,1,11,36,4,4,36,5,1,62,0,8,62,3,6,234,1,1,
/* out0115_em-eta15-phi5*/	13,42,4,4,70,0,10,70,2,1,70,3,5,48,1,5,48,2,1,36,5,11,37,5,4,62,3,1,38,4,4,38,5,5,234,0,1,234,1,7,
/* out0116_em-eta16-phi5*/	14,42,5,12,43,5,2,70,3,2,48,1,1,48,2,3,37,2,2,37,5,9,38,0,1,38,1,1,38,5,8,39,5,7,234,0,3,234,1,1,234,2,3,
/* out0117_em-eta17-phi5*/	15,28,0,1,28,2,4,43,2,1,43,5,11,44,1,1,17,3,1,37,2,5,38,0,6,222,2,1,234,0,1,234,2,4,39,2,4,39,5,6,40,0,2,40,1,1,
/* out0118_em-eta18-phi5*/	13,18,3,1,43,2,6,44,0,6,28,0,3,28,2,1,16,0,2,16,3,11,38,0,2,16,3,2,17,3,1,39,2,3,40,0,6,222,2,6,
/* out0119_em-eta19-phi5*/	10,18,0,1,18,3,11,19,3,1,44,0,3,16,0,6,16,0,4,16,3,9,40,0,1,222,0,2,222,2,1,
/* out0120_em-eta0-phi6*/	0,
/* out0121_em-eta1-phi6*/	0,
/* out0122_em-eta2-phi6*/	0,
/* out0123_em-eta3-phi6*/	0,
/* out0124_em-eta4-phi6*/	3,178,1,2,180,0,5,180,1,4,
/* out0125_em-eta5-phi6*/	5,160,1,5,162,0,3,180,0,11,180,1,5,180,2,15,
/* out0126_em-eta6-phi6*/	5,138,0,1,138,1,2,160,1,5,162,0,11,162,2,8,
/* out0127_em-eta7-phi6*/	4,138,1,13,138,2,1,140,0,5,162,2,2,
/* out0128_em-eta8-phi6*/	5,116,0,5,116,1,7,138,2,2,140,0,1,140,2,3,
/* out0129_em-eta9-phi6*/	3,116,1,7,116,2,7,86,4,5,
/* out0130_em-eta10-phi6*/	9,96,4,2,94,0,9,94,1,3,86,4,11,86,5,9,87,0,14,87,1,4,87,4,1,87,5,1,
/* out0131_em-eta11-phi6*/	12,96,4,14,96,5,9,97,0,11,97,1,4,94,0,1,94,1,1,94,2,9,86,2,2,87,2,5,87,3,6,87,4,15,87,5,4,
/* out0132_em-eta12-phi6*/	13,70,1,1,72,0,6,94,2,2,96,2,2,97,0,3,97,2,4,97,3,4,97,4,16,97,5,5,62,4,6,63,1,13,87,2,4,87,3,6,
/* out0133_em-eta13-phi6*/	11,70,4,6,71,1,10,97,2,5,97,3,7,72,0,4,72,2,3,62,1,2,62,2,10,63,0,10,63,1,1,63,4,1,
/* out0134_em-eta14-phi6*/	11,48,1,2,72,2,4,70,1,2,70,2,8,71,0,10,71,1,3,71,4,1,62,2,5,62,3,6,63,3,4,63,4,5,
/* out0135_em-eta15-phi6*/	12,48,1,3,50,0,2,70,2,7,70,3,5,71,3,3,71,4,5,37,5,1,38,1,1,39,1,5,62,3,3,63,3,6,234,1,6,
/* out0136_em-eta16-phi6*/	16,42,5,1,43,5,1,44,1,1,45,1,4,70,3,4,71,3,8,48,1,1,50,0,2,38,1,11,38,2,1,39,1,2,39,5,1,40,1,3,41,1,6,234,1,1,234,2,6,
/* out0137_em-eta17-phi6*/	16,28,0,3,50,2,1,44,1,10,44,2,1,45,1,3,38,0,4,38,1,3,38,2,3,38,3,1,222,0,1,222,2,2,234,2,3,236,0,1,40,1,11,40,2,2,41,1,1,
/* out0138_em-eta18-phi6*/	13,28,0,4,44,0,4,44,1,4,44,2,3,44,3,1,38,0,3,38,3,6,222,0,5,222,2,2,40,0,5,40,1,1,40,2,2,40,3,3,
/* out0139_em-eta19-phi6*/	9,18,0,15,44,0,3,44,3,12,16,0,3,38,3,3,16,0,11,40,0,2,40,3,7,222,0,2,
/* out0140_em-eta0-phi7*/	0,
/* out0141_em-eta1-phi7*/	0,
/* out0142_em-eta2-phi7*/	0,
/* out0143_em-eta3-phi7*/	0,
/* out0144_em-eta4-phi7*/	2,180,1,1,182,0,2,
/* out0145_em-eta5-phi7*/	6,162,0,1,162,1,2,180,1,6,180,2,1,182,0,13,182,2,8,
/* out0146_em-eta6-phi7*/	5,162,0,1,162,1,14,162,2,4,164,0,5,182,2,2,
/* out0147_em-eta7-phi7*/	4,140,0,10,140,1,8,162,2,2,164,2,1,
/* out0148_em-eta8-phi7*/	4,116,1,1,118,0,3,140,1,2,140,2,12,
/* out0149_em-eta9-phi7*/	3,116,1,1,118,0,11,118,2,4,
/* out0150_em-eta10-phi7*/	7,94,1,6,96,0,1,118,2,5,86,5,7,87,5,4,88,1,2,89,1,4,
/* out0151_em-eta11-phi7*/	11,96,5,7,97,5,2,98,1,1,99,1,4,94,1,6,94,2,2,96,0,3,87,2,6,87,5,7,88,0,8,88,1,13,
/* out0152_em-eta12-phi7*/	13,72,0,4,72,1,4,96,2,1,97,2,5,97,5,9,98,0,5,98,1,14,99,1,1,62,4,10,62,5,5,87,2,1,88,0,8,88,3,3,
/* out0153_em-eta13-phi7*/	12,70,4,10,70,5,3,97,2,2,98,0,11,98,3,3,72,0,1,72,1,4,72,2,2,62,5,7,63,0,6,63,4,5,63,5,5,
/* out0154_em-eta14-phi7*/	10,50,0,1,72,2,5,70,5,10,71,0,6,71,4,4,71,5,4,63,2,8,63,3,4,63,4,5,63,5,3,
/* out0155_em-eta15-phi7*/	10,50,0,5,71,2,6,71,3,3,71,4,6,71,5,4,38,4,6,39,1,5,63,2,3,63,3,2,236,1,1,
/* out0156_em-eta16-phi7*/	13,44,4,6,45,1,4,71,2,5,71,3,2,50,0,3,50,2,2,38,2,2,39,0,8,39,1,4,40,4,6,41,1,8,236,0,5,236,1,1,
/* out0157_em-eta17-phi7*/	11,44,2,1,45,0,7,45,1,5,50,2,3,38,2,8,39,0,1,39,4,2,40,2,3,41,0,9,41,1,1,236,0,5,
/* out0158_em-eta18-phi7*/	14,28,0,2,50,2,1,44,2,8,45,0,2,45,4,2,38,2,2,38,3,3,39,3,2,39,4,2,222,0,4,236,0,1,40,2,8,40,3,1,41,4,3,
/* out0159_em-eta19-phi7*/	11,44,2,3,44,3,3,45,3,11,45,4,2,38,3,3,39,3,5,222,0,1,40,2,1,40,3,5,41,3,4,41,4,1,
/* out0160_em-eta0-phi8*/	0,
/* out0161_em-eta1-phi8*/	0,
/* out0162_em-eta2-phi8*/	0,
/* out0163_em-eta3-phi8*/	0,
/* out0164_em-eta4-phi8*/	5,182,0,1,182,1,1,194,0,11,194,1,5,194,2,8,
/* out0165_em-eta5-phi8*/	7,182,1,15,182,2,5,184,0,8,184,2,2,194,0,4,194,1,8,194,2,4,
/* out0166_em-eta6-phi8*/	5,164,0,11,164,1,11,164,2,3,182,2,1,184,2,1,
/* out0167_em-eta7-phi8*/	3,140,1,4,142,0,7,164,2,11,
/* out0168_em-eta8-phi8*/	6,118,0,1,118,1,3,140,1,2,140,2,1,142,0,5,142,2,6,
/* out0169_em-eta9-phi8*/	3,118,0,1,118,1,12,118,2,2,
/* out0170_em-eta10-phi8*/	8,96,0,6,96,1,1,118,1,1,118,2,5,88,4,12,88,5,1,89,0,1,89,1,10,
/* out0171_em-eta11-phi8*/	10,98,4,12,99,1,7,96,0,6,96,1,1,96,2,4,88,1,1,88,2,13,89,0,13,89,1,2,89,4,5,
/* out0172_em-eta12-phi8*/	13,72,1,2,96,2,6,98,1,1,98,2,11,98,5,1,99,0,13,99,1,4,99,4,4,62,5,1,88,2,3,88,3,12,89,3,9,89,4,3,
/* out0173_em-eta13-phi8*/	12,72,1,5,74,0,3,98,2,5,98,3,11,99,3,7,99,4,4,62,5,3,63,5,7,64,1,8,65,1,4,88,3,1,89,3,1,
/* out0174_em-eta14-phi8*/	16,50,0,1,50,1,1,72,1,1,72,2,1,74,0,1,74,2,1,70,5,3,71,5,6,72,1,6,73,1,4,98,3,2,99,3,3,63,2,5,63,5,1,64,0,9,64,1,4,
/* out0175_em-eta15-phi8*/	11,50,0,2,50,1,4,71,2,4,71,5,2,72,0,8,72,1,6,38,4,10,38,5,1,64,0,5,40,4,1,236,1,4,
/* out0176_em-eta16-phi8*/	12,44,4,9,71,2,1,72,0,6,50,1,2,50,2,2,38,5,7,39,0,6,40,4,9,40,5,5,236,0,1,236,1,6,236,2,1,
/* out0177_em-eta17-phi8*/	12,44,4,1,44,5,7,45,0,5,50,2,4,39,0,1,39,4,10,39,5,1,40,5,3,41,0,7,41,4,3,236,0,2,236,2,3,
/* out0178_em-eta18-phi8*/	13,45,0,2,45,4,9,45,5,1,50,2,1,39,2,2,39,3,5,39,4,2,41,2,1,41,3,5,41,4,9,41,5,1,236,0,1,236,2,2,
/* out0179_em-eta19-phi8*/	7,45,2,2,45,3,5,45,4,3,39,2,1,39,3,4,41,2,2,41,3,7,
/* out0180_em-eta0-phi9*/	0,
/* out0181_em-eta1-phi9*/	0,
/* out0182_em-eta2-phi9*/	0,
/* out0183_em-eta3-phi9*/	0,
/* out0184_em-eta4-phi9*/	6,194,0,1,194,1,2,194,2,3,196,0,5,196,1,1,196,2,3,
/* out0185_em-eta5-phi9*/	8,184,0,8,184,1,16,184,2,6,194,1,1,194,2,1,196,0,7,196,1,7,196,2,1,
/* out0186_em-eta6-phi9*/	4,164,1,4,166,0,15,166,2,1,184,2,7,
/* out0187_em-eta7-phi9*/	6,142,0,3,142,1,9,164,1,1,164,2,1,166,0,1,166,2,7,
/* out0188_em-eta8-phi9*/	4,120,0,2,142,0,1,142,1,7,142,2,9,
/* out0189_em-eta9-phi9*/	3,120,0,13,120,2,1,142,2,1,
/* out0190_em-eta10-phi9*/	5,96,1,5,120,0,1,120,2,7,88,4,4,88,5,9,
/* out0191_em-eta11-phi9*/	9,98,4,4,98,5,6,96,1,9,96,2,1,88,5,6,89,0,2,89,2,3,89,4,7,89,5,16,
/* out0192_em-eta12-phi9*/	12,74,0,4,96,2,4,98,5,9,99,0,3,99,2,1,99,4,6,99,5,15,64,4,6,65,1,1,89,2,13,89,3,6,89,4,1,
/* out0193_em-eta13-phi9*/	11,72,4,4,99,2,15,99,3,6,99,4,2,99,5,1,74,0,7,64,1,2,64,2,1,64,4,2,65,0,7,65,1,11,
/* out0194_em-eta14-phi9*/	12,72,1,1,72,2,1,72,4,4,73,0,6,73,1,12,74,0,1,74,2,6,64,0,1,64,1,2,64,2,14,64,3,2,65,0,1,
/* out0195_em-eta15-phi9*/	12,50,1,4,74,2,1,72,0,1,72,1,3,72,2,14,72,3,1,73,0,2,38,5,1,64,0,1,64,2,1,64,3,13,236,1,1,
/* out0196_em-eta16-phi9*/	11,44,5,1,72,0,1,72,2,1,72,3,13,50,1,4,38,5,7,39,5,6,64,3,1,40,5,4,236,1,3,236,2,3,
/* out0197_em-eta17-phi9*/	10,44,5,8,45,5,5,72,3,2,50,1,1,50,2,2,39,2,3,39,5,9,40,5,4,41,5,9,236,2,6,
/* out0198_em-eta18-phi9*/	7,45,2,2,45,5,10,46,0,1,39,2,9,41,2,5,41,5,6,236,2,1,
/* out0199_em-eta19-phi9*/	4,45,2,12,46,0,1,39,2,1,41,2,8,
/* out0200_em-eta0-phi10*/	0,
/* out0201_em-eta1-phi10*/	0,
/* out0202_em-eta2-phi10*/	0,
/* out0203_em-eta3-phi10*/	0,
/* out0204_em-eta4-phi10*/	6,196,0,3,196,1,1,196,2,5,198,0,3,198,1,2,198,2,1,
/* out0205_em-eta5-phi10*/	8,186,0,16,186,1,8,186,2,6,196,0,1,196,1,7,196,2,7,198,0,1,198,1,1,
/* out0206_em-eta6-phi10*/	4,166,1,15,166,2,1,168,0,4,186,2,7,
/* out0207_em-eta7-phi10*/	6,144,0,9,144,1,3,166,1,1,166,2,7,168,0,1,168,2,1,
/* out0208_em-eta8-phi10*/	4,120,1,2,144,0,7,144,1,1,144,2,9,
/* out0209_em-eta9-phi10*/	3,120,1,13,120,2,1,144,2,1,
/* out0210_em-eta10-phi10*/	5,98,0,5,120,1,1,120,2,7,90,4,4,91,1,9,
/* out0211_em-eta11-phi10*/	9,100,4,4,101,1,6,98,0,9,98,2,1,90,0,3,90,1,16,90,2,7,91,0,2,91,1,6,
/* out0212_em-eta12-phi10*/	12,74,1,4,98,2,4,100,0,1,100,1,15,100,2,6,101,0,3,101,1,9,64,4,6,64,5,1,90,0,13,90,2,1,90,3,6,
/* out0213_em-eta13-phi10*/	11,72,4,4,100,0,15,100,1,1,100,2,2,100,3,6,74,1,7,64,4,2,64,5,11,65,0,7,65,4,1,65,5,2,
/* out0214_em-eta14-phi10*/	12,72,4,4,72,5,12,73,0,6,73,4,1,73,5,1,74,1,1,74,2,6,65,0,1,65,2,1,65,3,2,65,4,14,65,5,2,
/* out0215_em-eta15-phi10*/	12,52,0,4,74,2,1,73,0,2,73,2,1,73,3,1,73,4,14,73,5,2,41,1,1,65,2,1,65,3,13,65,4,1,238,1,1,
/* out0216_em-eta16-phi10*/	11,47,1,1,73,2,1,73,3,13,73,4,1,52,0,4,40,1,6,41,1,7,65,3,1,43,1,4,238,0,3,238,1,3,
/* out0217_em-eta17-phi10*/	10,46,1,5,47,1,8,73,3,2,52,0,1,52,2,2,40,0,3,40,1,9,42,1,9,43,1,4,238,0,6,
/* out0218_em-eta18-phi10*/	6,46,0,2,46,1,10,40,0,9,42,0,5,42,1,6,238,0,1,
/* out0219_em-eta19-phi10*/	3,46,0,10,40,0,1,42,0,8,
/* out0220_em-eta0-phi11*/	0,
/* out0221_em-eta1-phi11*/	0,
/* out0222_em-eta2-phi11*/	0,
/* out0223_em-eta3-phi11*/	0,
/* out0224_em-eta4-phi11*/	5,188,0,1,188,1,1,198,0,8,198,1,5,198,2,11,
/* out0225_em-eta5-phi11*/	7,186,1,8,186,2,2,188,0,15,188,2,5,198,0,4,198,1,8,198,2,4,
/* out0226_em-eta6-phi11*/	5,168,0,11,168,1,11,168,2,3,186,2,1,188,2,1,
/* out0227_em-eta7-phi11*/	3,144,1,7,146,0,4,168,2,11,
/* out0228_em-eta8-phi11*/	6,122,0,3,122,1,1,144,1,5,144,2,6,146,0,2,146,2,1,
/* out0229_em-eta9-phi11*/	3,122,0,12,122,1,1,122,2,2,
/* out0230_em-eta10-phi11*/	8,98,0,1,98,1,6,122,0,1,122,2,5,90,4,12,90,5,10,91,0,1,91,1,1,
/* out0231_em-eta11-phi11*/	10,100,4,12,100,5,7,98,0,1,98,1,6,98,2,4,90,2,5,90,5,2,91,0,13,91,4,13,91,5,1,
/* out0232_em-eta12-phi11*/	13,76,0,2,98,2,6,100,2,4,100,5,4,101,0,13,101,1,1,101,4,11,101,5,1,67,1,1,90,2,3,90,3,9,91,3,12,91,4,3,
/* out0233_em-eta13-phi11*/	12,74,1,3,76,0,5,100,2,4,100,3,7,101,3,11,101,4,5,64,5,4,65,5,8,66,1,7,67,1,3,90,3,1,91,3,1,
/* out0234_em-eta14-phi11*/	16,52,0,1,52,1,1,74,1,1,74,2,1,76,0,1,76,2,1,72,5,4,73,5,7,74,1,6,75,1,3,100,3,3,101,3,2,65,2,9,65,5,4,66,0,5,66,1,1,
/* out0235_em-eta15-phi11*/	11,52,0,4,52,1,2,73,2,8,73,5,6,74,0,4,74,1,2,40,4,10,41,1,1,65,2,5,42,4,1,238,1,4,
/* out0236_em-eta16-phi11*/	12,46,4,9,73,2,6,74,0,1,52,0,2,52,2,2,41,0,6,41,1,7,42,4,9,43,1,5,238,0,1,238,1,6,238,2,1,
/* out0237_em-eta17-phi11*/	12,46,4,1,47,0,5,47,1,7,52,2,4,40,1,1,40,2,10,41,0,1,42,2,3,43,0,7,43,1,3,238,0,3,238,2,2,
/* out0238_em-eta18-phi11*/	13,46,1,1,46,2,9,47,0,2,52,2,1,40,0,2,40,2,2,40,3,5,42,0,1,42,1,1,42,2,9,42,3,5,238,0,2,238,2,1,
/* out0239_em-eta19-phi11*/	7,46,0,2,46,2,3,46,3,5,40,0,1,40,3,4,42,0,2,42,3,7,
/* out0240_em-eta0-phi12*/	0,
/* out0241_em-eta1-phi12*/	0,
/* out0242_em-eta2-phi12*/	0,
/* out0243_em-eta3-phi12*/	0,
/* out0244_em-eta4-phi12*/	2,188,1,2,190,1,1,
/* out0245_em-eta5-phi12*/	7,170,0,2,170,1,1,188,1,13,188,2,8,190,0,13,190,1,1,190,2,1,
/* out0246_em-eta6-phi12*/	5,168,1,5,170,0,14,170,1,1,170,2,4,188,2,2,
/* out0247_em-eta7-phi12*/	4,146,0,8,146,1,10,168,2,1,170,2,2,
/* out0248_em-eta8-phi12*/	4,122,1,3,124,0,1,146,0,2,146,2,12,
/* out0249_em-eta9-phi12*/	3,122,1,11,122,2,4,124,0,1,
/* out0250_em-eta10-phi12*/	7,98,1,1,100,0,6,122,2,5,90,5,4,91,5,2,92,1,4,93,1,7,
/* out0251_em-eta11-phi12*/	11,100,5,4,101,5,1,102,1,2,103,1,7,98,1,3,100,0,6,100,2,2,91,2,8,91,5,13,92,0,6,92,1,7,
/* out0252_em-eta12-phi12*/	13,76,0,4,76,1,4,98,2,1,100,5,1,101,2,5,101,5,14,102,0,5,102,1,9,66,4,10,67,1,5,91,2,8,91,3,3,92,0,1,
/* out0253_em-eta13-phi12*/	12,74,4,10,75,1,3,101,2,11,101,3,3,102,0,2,76,0,4,76,1,1,76,2,2,66,1,5,66,2,5,67,0,6,67,1,7,
/* out0254_em-eta14-phi12*/	10,52,1,1,76,2,5,74,1,4,74,2,4,75,0,6,75,1,10,66,0,8,66,1,3,66,2,5,66,3,4,
/* out0255_em-eta15-phi12*/	10,52,1,5,74,0,6,74,1,4,74,2,6,74,3,3,40,4,6,40,5,5,66,0,3,66,3,2,238,1,1,
/* out0256_em-eta16-phi12*/	13,46,4,6,46,5,4,74,0,5,74,3,2,52,1,3,52,2,2,40,5,4,41,0,8,41,4,2,42,4,6,42,5,8,238,1,1,238,2,5,
/* out0257_em-eta17-phi12*/	11,46,5,5,47,0,7,47,4,1,52,2,3,40,2,2,41,0,1,41,4,8,42,5,1,43,0,9,43,4,3,238,2,5,
/* out0258_em-eta18-phi12*/	14,30,1,2,52,2,1,46,2,2,47,0,2,47,4,8,40,2,2,40,3,2,41,3,3,41,4,2,224,1,4,238,2,1,42,2,3,43,3,1,43,4,8,
/* out0259_em-eta19-phi12*/	11,46,2,2,46,3,11,47,3,3,47,4,3,40,3,5,41,3,3,224,1,1,42,2,1,42,3,4,43,3,5,43,4,1,
/* out0260_em-eta0-phi13*/	0,
/* out0261_em-eta1-phi13*/	0,
/* out0262_em-eta2-phi13*/	0,
/* out0263_em-eta3-phi13*/	0,
/* out0264_em-eta4-phi13*/	2,190,1,6,192,0,2,
/* out0265_em-eta5-phi13*/	5,170,1,3,172,0,5,190,0,3,190,1,8,190,2,15,
/* out0266_em-eta6-phi13*/	5,148,0,2,148,1,1,170,1,11,170,2,8,172,0,5,
/* out0267_em-eta7-phi13*/	4,146,1,5,148,0,13,148,2,1,170,2,2,
/* out0268_em-eta8-phi13*/	5,124,0,7,124,1,5,146,1,1,146,2,3,148,2,2,
/* out0269_em-eta9-phi13*/	3,124,0,7,124,2,7,92,4,5,
/* out0270_em-eta10-phi13*/	9,102,4,2,100,0,3,100,1,9,92,1,1,92,2,1,92,4,11,92,5,4,93,0,14,93,1,9,
/* out0271_em-eta11-phi13*/	12,102,4,14,102,5,4,103,0,11,103,1,9,100,0,1,100,1,1,100,2,9,92,0,5,92,1,4,92,2,15,92,3,6,93,4,2,
/* out0272_em-eta12-phi13*/	13,76,1,6,78,0,1,100,2,2,102,0,4,102,1,5,102,2,16,102,3,4,103,0,3,103,4,2,66,4,6,66,5,13,92,0,4,92,3,6,
/* out0273_em-eta13-phi13*/	11,74,4,6,74,5,10,102,0,5,102,3,7,76,1,4,76,2,3,66,2,1,66,5,1,67,0,10,67,4,10,67,5,2,
/* out0274_em-eta14-phi13*/	11,54,0,2,76,2,4,74,2,1,74,5,3,75,0,10,75,4,8,75,5,2,66,2,5,66,3,4,67,3,6,67,4,5,
/* out0275_em-eta15-phi13*/	11,52,1,2,54,0,3,74,2,5,74,3,3,75,3,5,75,4,7,40,5,5,41,5,1,42,1,1,66,3,6,67,3,3,
/* out0276_em-eta16-phi13*/	14,46,5,4,47,5,1,48,1,1,49,1,1,74,3,8,75,3,4,52,1,2,54,0,1,40,5,2,41,4,1,41,5,11,42,5,6,43,5,3,44,1,1,
/* out0277_em-eta17-phi13*/	15,30,1,3,52,2,1,46,5,3,47,4,1,47,5,10,41,2,4,41,3,1,41,4,3,41,5,3,224,1,1,224,2,2,238,2,1,42,5,1,43,4,2,43,5,11,
/* out0278_em-eta18-phi13*/	13,30,1,4,47,2,4,47,3,1,47,4,3,47,5,4,41,2,3,41,3,6,224,1,5,224,2,2,43,2,5,43,3,3,43,4,2,43,5,1,
/* out0279_em-eta19-phi13*/	9,20,4,15,47,2,3,47,3,12,18,4,3,41,3,3,18,4,11,43,2,2,43,3,7,224,1,2,
/* out0280_em-eta0-phi14*/	0,
/* out0281_em-eta1-phi14*/	0,
/* out0282_em-eta2-phi14*/	0,
/* out0283_em-eta3-phi14*/	0,
/* out0284_em-eta4-phi14*/	2,192,0,10,192,2,1,
/* out0285_em-eta5-phi14*/	5,172,0,4,172,1,14,174,0,1,192,0,4,192,2,13,
/* out0286_em-eta6-phi14*/	5,148,1,5,150,0,3,172,0,2,172,1,1,172,2,15,
/* out0287_em-eta7-phi14*/	5,126,0,1,148,0,1,148,1,10,148,2,9,150,0,1,
/* out0288_em-eta8-phi14*/	3,124,1,8,126,0,7,148,2,4,
/* out0289_em-eta9-phi14*/	5,102,0,4,124,1,3,124,2,8,126,0,1,92,5,1,
/* out0290_em-eta10-phi14*/	8,100,1,4,102,0,8,124,2,1,92,5,11,93,0,2,93,2,3,93,4,5,93,5,15,
/* out0291_em-eta11-phi14*/	17,78,0,3,78,1,1,100,1,2,100,2,3,102,2,1,102,5,12,103,0,2,103,2,2,103,4,3,103,5,14,68,4,1,69,1,1,92,3,1,93,2,9,93,3,12,93,4,9,93,5,1,
/* out0292_em-eta12-phi14*/	13,76,4,1,102,3,1,103,2,10,103,3,10,103,4,11,103,5,2,78,0,9,66,5,2,67,5,4,68,1,7,69,1,7,92,3,3,93,3,4,
/* out0293_em-eta13-phi14*/	16,54,1,1,76,1,1,76,2,1,78,0,2,78,2,2,74,5,3,75,5,3,76,1,6,77,1,8,102,3,4,103,3,6,67,2,8,67,4,1,67,5,10,68,0,2,68,1,2,
/* out0294_em-eta14-phi14*/	10,54,0,4,54,1,2,75,2,6,75,5,11,76,0,2,76,1,4,42,4,4,43,1,1,67,2,8,67,3,6,
/* out0295_em-eta15-phi14*/	11,48,4,4,75,2,10,75,3,5,75,4,1,54,0,5,54,2,1,42,1,4,43,1,11,67,3,1,44,4,4,45,1,5,
/* out0296_em-eta16-phi14*/	11,48,1,2,49,1,12,75,3,2,54,0,1,54,2,3,41,2,1,41,5,1,42,0,2,42,1,9,44,1,7,45,1,8,
/* out0297_em-eta17-phi14*/	13,30,1,1,30,2,4,47,5,1,48,0,1,48,1,11,19,5,1,41,2,6,42,0,5,224,2,1,43,2,2,43,5,1,44,0,4,44,1,6,
/* out0298_em-eta18-phi14*/	13,20,5,1,47,2,6,48,0,6,30,1,3,30,2,1,18,4,2,18,5,11,41,2,2,18,5,2,19,5,1,43,2,6,44,0,3,224,2,6,
/* out0299_em-eta19-phi14*/	10,20,4,1,20,5,11,21,5,1,47,2,3,18,4,6,18,4,4,18,5,9,43,2,1,224,1,2,224,2,1,
/* out0300_em-eta0-phi15*/	0,
/* out0301_em-eta1-phi15*/	0,
/* out0302_em-eta2-phi15*/	0,
/* out0303_em-eta3-phi15*/	0,
/* out0304_em-eta4-phi15*/	3,174,0,1,174,1,3,192,2,1,
/* out0305_em-eta5-phi15*/	4,174,0,14,174,1,9,174,2,9,192,2,1,
/* out0306_em-eta6-phi15*/	6,150,0,9,150,1,12,150,2,2,172,1,1,172,2,1,174,2,3,
/* out0307_em-eta7-phi15*/	4,126,0,1,126,1,7,150,0,3,150,2,10,
/* out0308_em-eta8-phi15*/	3,126,0,6,126,1,5,126,2,7,
/* out0309_em-eta9-phi15*/	3,102,0,1,102,1,9,126,2,5,
/* out0310_em-eta10-phi15*/	4,102,0,3,102,1,3,102,2,7,93,2,1,
/* out0311_em-eta11-phi15*/	7,78,1,7,102,2,4,68,4,15,68,5,4,69,0,1,69,1,2,93,2,3,
/* out0312_em-eta12-phi15*/	10,76,4,15,76,5,4,103,2,4,78,0,1,78,1,4,78,2,4,68,1,3,68,2,8,69,0,11,69,1,6,
/* out0313_em-eta13-phi15*/	10,54,1,1,78,2,6,76,1,2,76,2,6,77,0,12,77,1,8,68,0,12,68,1,4,68,2,4,68,3,4,
/* out0314_em-eta14-phi15*/	11,54,1,6,76,0,10,76,1,4,76,2,6,76,3,4,42,4,12,42,5,4,43,0,1,43,1,1,68,0,2,44,4,3,
/* out0315_em-eta15-phi15*/	12,48,4,12,48,5,4,76,0,4,54,1,2,54,2,3,42,2,3,43,0,11,43,1,3,44,4,9,44,5,4,45,0,3,45,1,2,
/* out0316_em-eta16-phi15*/	12,48,2,1,49,0,12,49,1,3,54,2,4,42,0,1,42,1,2,42,2,9,42,3,1,226,1,1,44,2,6,45,0,9,45,1,1,
/* out0317_em-eta17-phi15*/	14,30,2,4,54,2,1,48,0,1,48,1,2,48,2,11,19,5,2,42,0,8,42,3,3,226,0,1,226,1,3,44,0,3,44,1,2,44,2,6,44,3,3,
/* out0318_em-eta18-phi15*/	13,30,1,1,30,2,3,48,0,8,48,3,4,18,5,4,19,0,6,19,4,4,19,5,9,19,5,6,44,0,6,44,3,1,224,2,2,226,0,3,
/* out0319_em-eta19-phi15*/	17,20,5,4,21,0,16,21,4,12,21,5,11,30,1,1,18,4,5,18,5,1,19,0,6,19,1,2,18,4,1,18,5,5,19,0,15,19,1,16,19,4,4,19,5,5,224,1,1,224,2,2,
/* out0320_em-eta0-phi16*/	0,
/* out0321_em-eta1-phi16*/	0,
/* out0322_em-eta2-phi16*/	0,
/* out0323_em-eta3-phi16*/	0,
/* out0324_em-eta4-phi16*/	1,176,0,7,
/* out0325_em-eta5-phi16*/	6,152,0,5,152,1,7,174,1,4,174,2,4,176,0,8,176,2,8,
/* out0326_em-eta6-phi16*/	6,128,1,2,150,1,4,150,2,1,152,0,11,152,1,1,152,2,7,
/* out0327_em-eta7-phi16*/	5,126,1,1,128,0,14,128,1,4,128,2,1,150,2,3,
/* out0328_em-eta8-phi16*/	6,104,0,4,104,1,3,126,1,3,126,2,4,128,0,2,128,2,3,
/* out0329_em-eta9-phi16*/	3,102,1,2,104,0,11,104,2,1,
/* out0330_em-eta10-phi16*/	7,80,0,4,80,1,1,102,1,2,102,2,4,104,0,1,104,2,1,71,1,1,
/* out0331_em-eta11-phi16*/	7,78,1,1,80,0,9,68,5,12,69,0,1,69,5,10,70,1,2,71,1,2,
/* out0332_em-eta12-phi16*/	15,56,0,1,78,1,3,78,2,2,80,0,1,80,2,1,76,5,12,77,5,7,78,1,2,79,1,2,68,2,1,69,0,3,69,2,2,69,3,3,69,4,15,69,5,5,
/* out0333_em-eta13-phi16*/	12,56,0,6,78,2,2,76,2,1,77,0,4,77,2,1,77,3,2,77,4,14,77,5,7,68,2,3,68,3,10,69,3,9,69,4,1,
/* out0334_em-eta14-phi16*/	11,54,1,2,56,0,4,76,2,3,76,3,8,77,3,10,77,4,2,42,5,12,43,0,1,43,5,5,68,3,2,44,5,3,
/* out0335_em-eta15-phi16*/	13,32,0,1,54,1,2,54,2,2,48,5,12,49,5,4,76,3,4,43,0,3,43,4,10,43,5,2,44,5,9,45,0,2,45,4,1,45,5,6,
/* out0336_em-eta16-phi16*/	14,32,0,3,54,2,2,49,0,4,49,4,9,49,5,3,42,2,4,42,3,1,43,3,3,43,4,6,226,1,4,44,2,1,45,0,2,45,4,12,45,5,1,
/* out0337_em-eta17-phi16*/	14,30,2,1,32,0,3,48,2,4,49,3,3,49,4,7,19,2,1,42,3,10,43,3,1,226,0,1,226,1,5,44,2,3,44,3,4,45,3,3,45,4,3,
/* out0338_em-eta18-phi16*/	11,30,2,3,48,3,11,49,3,1,19,2,7,19,3,1,19,4,6,19,5,4,19,2,5,19,5,1,44,3,7,226,0,5,
/* out0339_em-eta19-phi16*/	16,21,2,8,21,3,1,21,4,4,21,5,4,30,1,1,18,1,4,18,3,4,19,0,4,19,1,8,19,4,5,19,0,1,19,2,3,19,3,5,19,4,11,19,5,3,226,0,2,
/* out0340_em-eta0-phi17*/	0,
/* out0341_em-eta1-phi17*/	0,
/* out0342_em-eta2-phi17*/	0,
/* out0343_em-eta3-phi17*/	0,
/* out0344_em-eta4-phi17*/	4,154,0,1,154,1,4,176,0,1,176,2,3,
/* out0345_em-eta5-phi17*/	5,152,1,7,154,0,15,154,1,3,154,2,4,176,2,5,
/* out0346_em-eta6-phi17*/	5,128,1,2,130,0,12,130,1,2,152,1,1,152,2,9,
/* out0347_em-eta7-phi17*/	4,106,0,3,128,1,8,128,2,8,130,0,3,
/* out0348_em-eta8-phi17*/	3,104,1,9,106,0,5,128,2,4,
/* out0349_em-eta9-phi17*/	3,104,1,4,104,2,11,70,4,1,
/* out0350_em-eta10-phi17*/	7,80,1,10,82,0,1,104,2,2,70,4,15,70,5,3,71,0,7,71,1,10,
/* out0351_em-eta11-phi17*/	13,78,4,16,78,5,4,79,0,5,79,1,8,80,0,2,80,1,2,80,2,6,69,5,1,70,0,5,70,1,14,70,2,7,71,0,2,71,1,3,
/* out0352_em-eta12-phi17*/	11,56,1,5,80,2,4,77,5,1,78,0,2,78,1,14,78,2,7,79,0,4,79,1,6,44,4,7,69,2,13,70,0,7,
/* out0353_em-eta13-phi17*/	12,50,4,5,77,2,13,77,5,1,78,0,10,56,0,3,56,1,4,56,2,1,44,4,3,45,0,1,45,1,15,69,2,1,69,3,4,
/* out0354_em-eta14-phi17*/	9,50,4,5,51,1,13,77,2,2,77,3,4,56,0,2,56,2,4,43,5,5,44,0,2,44,1,13,
/* out0355_em-eta15-phi17*/	13,32,0,1,32,1,3,56,2,1,49,5,4,50,0,1,50,1,13,51,1,2,43,2,11,43,5,4,44,0,1,228,1,1,45,2,2,45,5,7,
/* out0356_em-eta16-phi17*/	15,32,0,3,32,1,1,49,2,10,49,5,5,50,0,2,20,4,1,21,1,1,43,2,4,43,3,8,226,1,2,226,2,2,228,0,1,45,2,11,45,3,2,45,5,2,
/* out0357_em-eta17-phi17*/	15,22,4,1,49,2,5,49,3,7,32,0,3,19,2,1,20,1,1,21,1,5,42,3,1,43,3,4,20,4,1,21,1,2,45,2,2,45,3,9,226,1,1,226,2,5,
/* out0358_em-eta18-phi17*/	15,23,1,5,48,3,1,49,3,5,32,0,2,32,2,1,19,2,7,19,3,5,20,1,2,19,2,3,20,1,3,21,1,4,44,3,1,45,3,2,226,0,2,226,2,3,
/* out0359_em-eta19-phi17*/	13,21,2,8,21,3,14,22,1,3,18,1,10,18,3,10,19,1,5,19,3,6,19,4,1,19,2,5,19,3,9,19,4,1,20,1,1,226,0,2,
/* out0360_em-eta0-phi18*/	0,
/* out0361_em-eta1-phi18*/	0,
/* out0362_em-eta2-phi18*/	0,
/* out0363_em-eta3-phi18*/	0,
/* out0364_em-eta4-phi18*/	4,154,1,4,156,0,12,156,1,6,156,2,7,
/* out0365_em-eta5-phi18*/	8,130,1,1,132,0,10,132,1,2,154,1,5,154,2,12,156,0,2,156,1,7,156,2,5,
/* out0366_em-eta6-phi18*/	5,108,0,1,130,0,1,130,1,13,130,2,9,132,0,3,
/* out0367_em-eta7-phi18*/	4,106,0,1,106,1,12,108,0,2,130,2,7,
/* out0368_em-eta8-phi18*/	3,106,0,7,106,1,1,106,2,10,
/* out0369_em-eta9-phi18*/	6,82,0,7,82,1,7,104,2,1,106,2,1,70,5,4,71,5,1,
/* out0370_em-eta10-phi18*/	10,78,5,1,79,5,1,80,1,2,82,0,8,82,2,3,70,5,9,71,0,6,71,2,1,71,4,8,71,5,15,
/* out0371_em-eta11-phi18*/	14,58,0,4,58,1,1,80,1,1,80,2,4,78,5,11,79,0,6,79,2,1,79,4,6,79,5,15,70,2,9,70,3,9,71,0,1,71,3,7,71,4,8,
/* out0372_em-eta12-phi18*/	12,56,1,3,58,0,5,80,2,1,78,2,9,78,3,6,79,0,1,79,3,7,79,4,10,44,4,5,44,5,13,70,0,4,70,3,6,
/* out0373_em-eta13-phi18*/	12,50,4,5,50,5,11,78,0,4,78,3,9,56,1,4,56,2,3,44,2,3,44,4,1,44,5,1,45,0,15,45,1,1,45,4,3,
/* out0374_em-eta14-phi18*/	12,50,2,1,50,4,1,50,5,3,51,0,16,51,1,1,51,4,2,56,2,6,44,0,4,44,1,3,44,2,10,44,3,3,228,1,2,
/* out0375_em-eta15-phi18*/	10,32,1,4,56,2,1,50,0,2,50,1,3,50,2,12,50,3,2,20,4,6,43,2,1,44,0,9,228,1,8,
/* out0376_em-eta16-phi18*/	13,22,4,5,49,2,1,50,0,11,50,3,1,32,1,4,32,2,1,20,4,8,21,0,1,21,1,5,20,4,10,45,2,1,228,0,6,228,1,1,
/* out0377_em-eta17-phi18*/	14,22,4,9,23,0,1,23,1,4,32,2,3,20,1,3,20,2,1,21,0,2,21,1,5,20,4,4,21,0,2,21,1,7,214,1,1,226,2,4,228,0,1,
/* out0378_em-eta18-phi18*/	13,22,1,2,22,2,1,23,0,2,23,1,7,32,2,3,20,0,1,20,1,8,20,1,5,20,2,1,21,0,1,21,1,3,214,1,2,226,2,2,
/* out0379_em-eta19-phi18*/	12,21,3,1,22,0,14,22,1,9,18,1,2,18,3,2,19,1,1,19,3,4,20,0,3,19,3,2,20,0,3,20,1,5,214,1,2,
/* out0380_em-eta0-phi19*/	0,
/* out0381_em-eta1-phi19*/	0,
/* out0382_em-eta2-phi19*/	0,
/* out0383_em-eta3-phi19*/	0,
/* out0384_em-eta4-phi19*/	3,134,1,9,156,0,2,156,2,2,
/* out0385_em-eta5-phi19*/	9,110,0,1,132,0,2,132,1,14,132,2,9,134,0,16,134,1,1,134,2,1,156,1,3,156,2,2,
/* out0386_em-eta6-phi19*/	5,108,0,4,108,1,13,110,0,1,132,0,1,132,2,7,
/* out0387_em-eta7-phi19*/	4,84,1,2,106,1,3,108,0,9,108,2,8,
/* out0388_em-eta8-phi19*/	3,84,0,10,84,1,2,106,2,5,
/* out0389_em-eta9-phi19*/	3,82,1,9,82,2,3,84,0,3,
/* out0390_em-eta10-phi19*/	5,58,1,2,60,0,1,82,2,10,46,4,6,71,2,11,
/* out0391_em-eta11-phi19*/	8,52,4,5,79,2,9,58,0,2,58,1,9,46,4,6,47,1,14,71,2,4,71,3,9,
/* out0392_em-eta12-phi19*/	13,52,4,8,53,1,12,79,2,6,79,3,8,58,0,4,58,2,5,44,5,2,45,2,1,45,5,12,46,0,1,46,1,10,47,1,1,70,3,1,
/* out0393_em-eta13-phi19*/	17,34,0,2,34,1,3,58,0,1,58,2,2,50,5,2,51,2,1,51,5,10,52,0,1,52,1,10,53,1,3,78,3,1,79,3,1,45,2,5,45,3,3,45,4,11,45,5,4,230,1,2,
/* out0394_em-eta14-phi19*/	13,34,0,6,51,2,5,51,3,2,51,4,10,51,5,6,44,2,3,44,3,8,45,3,7,45,4,2,228,1,2,228,2,2,230,0,1,230,1,2,
/* out0395_em-eta15-phi19*/	11,32,1,1,34,0,4,50,2,3,50,3,6,51,3,8,51,4,4,20,4,1,20,5,10,44,3,5,228,1,2,228,2,5,
/* out0396_em-eta16-phi19*/	11,22,4,1,22,5,8,50,3,7,32,1,3,32,2,2,20,5,4,21,0,9,20,4,1,20,5,13,228,0,5,228,2,2,
/* out0397_em-eta17-phi19*/	11,22,5,6,23,0,8,32,2,4,20,2,7,21,0,4,21,4,1,20,5,1,21,0,11,21,4,1,214,2,4,228,0,2,
/* out0398_em-eta18-phi19*/	12,22,2,6,23,0,5,23,4,1,32,2,2,20,0,3,20,1,2,20,2,4,20,3,1,20,2,9,21,0,2,214,1,3,214,2,1,
/* out0399_em-eta19-phi19*/	10,22,0,2,22,1,2,22,2,5,22,3,2,20,0,7,20,0,5,20,1,2,20,2,2,20,3,1,214,1,3,
/* out0400_em-eta0-phi20*/	0,
/* out0401_em-eta1-phi20*/	0,
/* out0402_em-eta2-phi20*/	0,
/* out0403_em-eta3-phi20*/	0,
/* out0404_em-eta4-phi20*/	3,112,1,2,134,1,6,134,2,2,
/* out0405_em-eta5-phi20*/	6,110,0,5,110,1,14,110,2,2,112,0,5,112,1,4,134,2,13,
/* out0406_em-eta6-phi20*/	6,86,0,1,86,1,4,108,1,3,108,2,2,110,0,9,110,2,8,
/* out0407_em-eta7-phi20*/	3,84,1,4,86,0,11,108,2,6,
/* out0408_em-eta8-phi20*/	3,84,0,2,84,1,8,84,2,9,
/* out0409_em-eta9-phi20*/	4,60,0,2,60,1,7,84,0,1,84,2,6,
/* out0410_em-eta10-phi20*/	6,60,0,11,60,1,1,60,2,1,46,4,3,46,5,15,47,5,5,
/* out0411_em-eta11-phi20*/	14,36,0,1,58,1,4,58,2,3,60,0,2,60,2,1,52,4,2,52,5,13,53,5,5,46,2,8,46,4,1,46,5,1,47,0,16,47,1,1,47,4,7,
/* out0412_em-eta12-phi20*/	15,36,0,2,58,2,6,52,2,4,52,4,1,52,5,3,53,0,16,53,1,1,53,4,7,53,5,1,45,2,1,46,0,12,46,1,6,46,2,7,46,3,3,230,1,1,
/* out0413_em-eta13-phi20*/	12,34,1,7,52,0,10,52,1,6,52,2,10,52,3,3,22,4,11,23,1,1,45,2,9,46,0,2,22,4,2,230,1,10,230,2,1,
/* out0414_em-eta14-phi20*/	13,24,4,10,51,2,9,52,0,4,34,0,2,34,1,2,34,2,2,22,1,2,23,1,12,45,3,6,22,4,9,23,1,4,230,0,8,230,1,1,
/* out0415_em-eta15-phi20*/	16,24,1,1,24,4,1,25,1,12,51,2,1,51,3,6,34,0,2,34,2,3,20,5,2,21,5,9,22,1,5,21,5,1,22,1,4,23,1,9,216,1,2,228,2,4,230,0,2,
/* out0416_em-eta16-phi20*/	15,14,1,1,14,2,1,34,2,1,22,5,2,23,5,8,24,1,6,25,1,1,21,4,7,21,5,7,20,5,2,21,5,12,22,1,2,216,1,3,228,0,1,228,2,3,
/* out0417_em-eta17-phi20*/	10,14,1,3,23,4,6,23,5,8,20,2,2,21,3,1,21,4,8,21,4,10,21,5,3,214,2,5,216,0,1,
/* out0418_em-eta18-phi20*/	14,14,1,2,22,2,1,23,3,1,23,4,9,20,2,2,20,3,7,21,3,1,20,2,4,20,3,1,21,3,1,21,4,5,214,0,2,214,1,1,214,2,3,
/* out0419_em-eta19-phi20*/	8,22,2,3,22,3,7,23,3,1,20,0,2,20,3,3,20,0,8,20,3,9,214,1,3,
/* out0420_em-eta0-phi21*/	0,
/* out0421_em-eta1-phi21*/	0,
/* out0422_em-eta2-phi21*/	0,
/* out0423_em-eta3-phi21*/	0,
/* out0424_em-eta4-phi21*/	1,112,1,4,
/* out0425_em-eta5-phi21*/	7,88,0,4,88,1,8,110,1,2,110,2,3,112,0,11,112,1,6,112,2,16,
/* out0426_em-eta6-phi21*/	4,86,1,10,86,2,1,88,0,12,110,2,3,
/* out0427_em-eta7-phi21*/	4,62,1,1,86,0,3,86,1,2,86,2,15,
/* out0428_em-eta8-phi21*/	4,62,0,9,62,1,7,84,2,1,86,0,1,
/* out0429_em-eta9-phi21*/	3,60,1,7,60,2,1,62,0,7,
/* out0430_em-eta10-phi21*/	4,60,1,1,60,2,11,47,2,5,47,5,8,
/* out0431_em-eta11-phi21*/	11,36,0,1,36,1,7,60,2,2,53,2,3,53,5,6,47,2,11,47,3,11,47,4,9,47,5,3,232,0,3,232,1,3,
/* out0432_em-eta12-phi21*/	16,36,0,8,36,1,1,53,2,13,53,3,8,53,4,8,53,5,4,22,4,1,22,5,6,46,0,1,46,2,1,46,3,13,47,3,5,230,2,1,232,0,13,232,1,1,232,2,7,
/* out0433_em-eta13-phi21*/	16,24,5,4,52,0,1,52,2,2,52,3,13,53,3,8,53,4,1,34,1,4,36,0,4,22,4,4,22,5,10,23,0,9,23,1,1,22,4,2,22,5,11,230,2,10,232,2,1,
/* out0434_em-eta14-phi21*/	15,24,4,5,24,5,12,25,0,7,34,2,6,22,1,2,22,2,7,23,0,7,23,1,2,22,4,3,22,5,5,23,0,13,23,1,2,216,1,1,230,0,5,230,2,4,
/* out0435_em-eta15-phi21*/	15,14,2,1,34,2,4,24,1,1,24,2,7,25,0,9,25,1,3,21,2,1,22,0,7,22,1,7,22,2,1,22,1,6,22,2,8,23,0,3,23,1,1,216,1,7,
/* out0436_em-eta16-phi21*/	11,14,2,5,24,0,6,24,1,8,24,2,1,21,2,13,22,0,1,21,2,4,22,0,8,22,1,4,216,0,3,216,1,3,
/* out0437_em-eta17-phi21*/	9,14,1,3,23,2,12,24,0,2,21,2,2,21,3,9,21,2,12,21,3,2,214,2,2,216,0,4,
/* out0438_em-eta18-phi21*/	8,14,1,2,23,2,4,23,3,8,20,3,4,21,3,5,21,3,10,214,0,8,214,2,1,
/* out0439_em-eta19-phi21*/	7,22,3,4,23,3,6,20,3,1,20,3,5,21,3,3,214,0,6,214,1,1,
/* out0440_em-eta0-phi22*/	0,
/* out0441_em-eta1-phi22*/	0,
/* out0442_em-eta2-phi22*/	0,
/* out0443_em-eta3-phi22*/	0,
/* out0444_em-eta4-phi22*/	1,90,1,5,
/* out0445_em-eta5-phi22*/	7,66,0,3,66,1,2,88,1,8,88,2,4,90,0,16,90,1,10,90,2,9,
/* out0446_em-eta6-phi22*/	4,64,0,1,64,1,10,66,0,3,88,2,12,
/* out0447_em-eta7-phi22*/	4,62,1,1,64,0,15,64,1,2,64,2,3,
/* out0448_em-eta8-phi22*/	4,40,0,1,62,1,7,62,2,9,64,2,1,
/* out0449_em-eta9-phi22*/	3,38,0,1,38,1,7,62,2,7,
/* out0450_em-eta10-phi22*/	4,38,0,11,38,1,1,24,4,5,24,5,8,
/* out0451_em-eta11-phi22*/	14,26,4,3,26,5,6,36,1,7,36,2,1,38,0,2,24,4,11,24,5,3,25,0,9,25,1,11,24,4,11,24,5,10,25,0,1,220,0,1,232,1,5,
/* out0452_em-eta12-phi22*/	20,26,4,13,26,5,4,27,0,8,27,1,8,36,1,1,36,2,8,23,2,1,23,5,6,24,0,1,24,1,13,24,2,1,25,1,5,218,1,1,232,1,7,232,2,6,24,1,2,24,2,2,24,4,5,25,0,8,25,1,15,
/* out0453_em-eta13-phi22*/	19,16,1,4,36,2,4,25,5,4,26,0,1,26,1,13,26,2,2,27,0,1,27,1,8,23,2,4,23,3,1,23,4,9,23,5,10,23,2,2,23,5,11,24,0,1,24,1,11,25,1,1,218,1,10,232,2,2,
/* out0454_em-eta14-phi22*/	15,16,0,6,25,2,5,25,4,7,25,5,12,22,2,7,22,3,2,23,3,2,23,4,7,23,2,3,23,3,2,23,4,13,23,5,5,216,2,1,218,0,5,218,1,4,
/* out0455_em-eta15-phi22*/	15,14,2,1,16,0,4,24,2,7,24,3,1,25,3,3,25,4,9,0,4,1,22,0,7,22,2,1,22,3,7,22,2,8,22,3,6,23,3,1,23,4,3,216,2,7,
/* out0456_em-eta16-phi22*/	11,14,2,5,24,0,6,24,2,1,24,3,8,0,4,13,22,0,1,0,4,4,22,0,8,22,3,4,216,0,3,216,2,3,
/* out0457_em-eta17-phi22*/	11,0,4,12,24,0,2,14,0,3,14,1,2,14,2,1,0,4,2,1,1,9,0,4,12,1,1,2,206,2,2,216,0,4,
/* out0458_em-eta18-phi22*/	8,0,4,4,1,1,8,14,1,2,0,1,4,1,1,5,1,1,10,206,1,3,206,2,1,
/* out0459_em-eta19-phi22*/	7,0,1,4,1,1,6,22,3,3,0,1,1,0,1,5,1,1,3,206,1,3,
/* out0460_em-eta0-phi23*/	0,
/* out0461_em-eta1-phi23*/	0,
/* out0462_em-eta2-phi23*/	0,
/* out0463_em-eta3-phi23*/	0,
/* out0464_em-eta4-phi23*/	3,68,1,8,90,1,1,90,2,1,
/* out0465_em-eta5-phi23*/	7,66,0,2,66,1,14,66,2,5,68,0,16,68,1,5,68,2,2,90,2,6,
/* out0466_em-eta6-phi23*/	6,42,0,2,42,1,3,64,1,4,64,2,1,66,0,8,66,2,9,
/* out0467_em-eta7-phi23*/	3,40,1,4,42,0,6,64,2,11,
/* out0468_em-eta8-phi23*/	3,40,0,9,40,1,8,40,2,2,
/* out0469_em-eta9-phi23*/	4,38,1,7,38,2,2,40,0,6,40,2,1,
/* out0470_em-eta10-phi23*/	6,38,0,1,38,1,1,38,2,11,24,5,5,25,2,3,25,5,15,
/* out0471_em-eta11-phi23*/	21,18,0,3,18,1,4,36,2,1,38,0,1,38,2,2,26,5,5,27,2,2,27,5,13,24,2,8,25,0,7,25,2,1,25,3,1,25,4,16,25,5,1,24,5,6,25,0,2,25,2,4,25,4,5,25,5,16,220,0,3,220,1,5,
/* out0472_em-eta12-phi23*/	23,18,0,6,36,2,2,26,2,4,26,5,1,27,0,7,27,2,1,27,3,1,27,4,16,27,5,3,2,4,1,24,0,12,24,1,3,24,2,7,24,3,6,218,2,1,220,0,12,220,1,1,220,2,7,24,2,13,24,3,2,25,0,5,25,3,1,25,4,11,
/* out0473_em-eta13-phi23*/	17,16,1,7,26,0,10,26,1,3,26,2,10,26,3,6,2,4,9,23,2,11,23,3,1,24,0,2,2,4,3,23,2,2,24,0,14,24,1,3,24,2,1,24,3,4,218,1,1,218,2,10,
/* out0474_em-eta14-phi23*/	15,2,4,9,25,2,10,26,0,4,16,0,2,16,1,2,16,2,2,3,1,6,22,3,2,23,3,12,2,4,7,3,1,2,23,2,9,23,3,4,218,0,8,218,2,1,
/* out0475_em-eta15-phi23*/	17,2,4,1,3,1,6,24,3,1,25,2,1,25,3,12,16,0,3,16,2,2,0,5,9,1,5,2,22,3,5,0,5,1,3,1,4,22,3,4,23,3,9,208,1,4,216,2,2,218,0,2,
/* out0476_em-eta16-phi23*/	15,0,5,8,1,5,2,24,3,6,25,3,1,14,0,3,14,2,2,16,0,1,0,5,7,1,0,7,0,5,12,1,5,2,22,3,2,208,0,1,208,1,3,216,2,3,
/* out0477_em-eta17-phi23*/	10,0,5,8,1,0,6,14,0,8,0,2,2,1,0,8,1,1,1,0,5,3,1,0,10,206,2,5,216,0,1,
/* out0478_em-eta18-phi23*/	14,0,2,1,1,0,9,1,1,1,14,0,1,14,1,1,0,1,7,0,2,2,1,1,1,0,1,1,0,2,4,1,0,5,1,1,1,206,1,2,206,2,3,
/* out0479_em-eta19-phi23*/	8,0,1,7,0,2,3,1,1,1,0,0,2,0,1,3,0,0,8,0,1,9,206,1,3,
/* out0480_em-eta0-phi24*/	0,
/* out0481_em-eta1-phi24*/	0,
/* out0482_em-eta2-phi24*/	0,
/* out0483_em-eta3-phi24*/	0,
/* out0484_em-eta4-phi24*/	4,46,0,2,46,2,2,68,1,3,68,2,6,
/* out0485_em-eta5-phi24*/	7,44,0,9,44,1,14,44,2,2,46,0,2,46,1,3,66,2,1,68,2,8,
/* out0486_em-eta6-phi24*/	5,42,1,13,42,2,4,44,0,7,44,2,1,66,2,1,
/* out0487_em-eta7-phi24*/	4,22,1,3,40,1,2,42,0,8,42,2,9,
/* out0488_em-eta8-phi24*/	3,22,0,5,40,1,2,40,2,10,
/* out0489_em-eta9-phi24*/	3,20,0,3,20,1,9,40,2,3,
/* out0490_em-eta10-phi24*/	5,18,1,2,20,0,10,38,2,1,4,4,11,25,2,6,
/* out0491_em-eta11-phi24*/	13,4,4,9,27,2,5,18,1,9,18,2,2,4,4,4,5,1,9,25,2,6,25,3,14,4,4,14,5,1,1,25,2,11,212,0,2,220,1,7,
/* out0492_em-eta12-phi24*/	23,4,4,6,5,1,8,27,2,8,27,3,12,18,0,5,18,2,4,2,4,1,2,5,12,3,5,2,4,1,1,24,0,1,24,3,10,25,3,1,3,5,1,4,1,1,4,4,1,5,1,8,24,3,5,25,2,1,25,3,15,210,1,2,220,1,3,220,2,8,
/* out0493_em-eta13-phi24*/	25,2,4,1,2,5,10,3,5,2,4,1,1,5,1,1,26,0,1,26,3,10,27,3,3,16,1,3,16,2,2,18,0,2,18,2,1,2,4,5,2,5,4,3,0,11,3,1,3,2,4,3,2,5,15,3,0,2,3,5,2,24,0,1,24,3,5,210,1,8,218,2,2,220,2,1,
/* out0494_em-eta14-phi24*/	20,2,4,5,2,5,6,3,0,10,3,1,2,16,2,6,2,1,8,2,2,3,3,0,2,3,1,7,2,2,1,2,4,3,2,5,1,3,0,12,3,1,6,208,1,2,208,2,2,210,0,2,210,1,2,218,0,1,218,2,2,
/* out0495_em-eta15-phi24*/	14,0,1,1,16,2,4,2,1,6,2,2,3,3,0,4,3,1,8,1,2,1,1,5,10,2,1,5,2,1,12,2,2,2,3,1,4,208,1,5,208,2,2,
/* out0496_em-eta16-phi24*/	12,1,2,1,1,5,8,2,1,7,0,0,2,0,1,3,1,4,9,1,5,4,1,2,1,1,5,13,2,1,1,208,0,5,208,1,2,
/* out0497_em-eta17-phi24*/	11,1,4,8,1,5,6,0,0,4,0,2,7,1,0,1,1,4,4,1,0,1,1,4,11,1,5,1,206,2,4,208,0,2,
/* out0498_em-eta18-phi24*/	14,0,2,6,1,0,1,1,4,5,0,0,2,14,0,1,0,0,3,0,1,1,0,2,4,0,3,2,0,2,9,1,4,2,206,0,7,206,1,1,206,2,1,
/* out0499_em-eta19-phi24*/	10,0,0,2,0,1,5,0,2,5,0,3,2,0,0,7,0,0,5,0,1,1,0,2,2,0,3,2,206,1,3,
/* out0500_em-eta0-phi25*/	0,
/* out0501_em-eta1-phi25*/	0,
/* out0502_em-eta2-phi25*/	0,
/* out0503_em-eta3-phi25*/	0,
/* out0504_em-eta4-phi25*/	4,26,1,4,46,0,7,46,1,6,46,2,12,
/* out0505_em-eta5-phi25*/	8,24,1,1,26,0,12,26,1,5,44,1,2,44,2,10,46,0,5,46,1,7,46,2,2,
/* out0506_em-eta6-phi25*/	5,24,0,9,24,1,13,24,2,1,42,2,1,44,2,3,
/* out0507_em-eta7-phi25*/	4,22,1,12,22,2,1,24,0,7,42,2,2,
/* out0508_em-eta8-phi25*/	3,22,0,10,22,1,1,22,2,7,
/* out0509_em-eta9-phi25*/	6,6,0,1,20,1,7,20,2,7,22,0,1,4,5,1,5,5,4,
/* out0510_em-eta10-phi25*/	12,4,1,2,20,0,3,20,2,8,4,5,1,5,5,1,4,4,1,4,5,15,5,0,8,5,4,6,5,5,9,4,5,6,5,5,9,
/* out0511_em-eta11-phi25*/	23,4,0,4,4,1,1,18,1,1,18,2,4,4,4,1,4,5,15,5,0,6,5,4,6,5,5,11,4,1,9,4,2,9,5,0,8,5,1,7,5,4,1,4,2,2,4,4,1,4,5,10,5,0,14,5,1,2,5,4,7,5,5,3,212,0,10,212,2,1,
/* out0512_em-eta12-phi25*/	21,2,1,3,4,0,1,18,2,5,4,1,6,4,2,9,5,0,10,5,1,7,5,4,1,3,2,5,3,5,13,4,0,4,4,1,6,4,0,2,4,1,15,4,2,7,5,0,2,5,1,5,210,1,1,210,2,6,212,0,2,212,2,7,
/* out0513_em-eta13-phi25*/	19,2,0,3,2,1,4,3,2,5,3,5,11,4,0,4,4,1,9,2,2,3,3,0,3,3,2,1,3,3,1,3,4,15,3,5,1,3,2,6,3,4,5,3,5,13,4,0,1,210,0,4,210,1,3,210,2,5,
/* out0514_em-eta14-phi25*/	17,2,0,6,2,2,1,3,0,2,3,2,1,3,3,1,3,4,16,3,5,3,2,0,4,2,1,3,2,2,10,2,3,3,2,2,8,3,0,2,3,3,1,3,4,11,208,2,2,210,0,7,
/* out0515_em-eta15-phi25*/	13,0,1,4,2,0,1,2,0,2,2,1,2,2,2,12,2,3,3,1,2,6,2,0,9,2,0,8,2,1,3,2,2,5,2,3,3,208,2,8,
/* out0516_em-eta16-phi25*/	12,1,2,5,2,0,11,2,1,1,0,0,1,0,1,4,1,2,8,1,3,5,1,4,1,1,2,10,2,0,5,208,0,6,208,2,1,
/* out0517_em-eta17-phi25*/	14,1,2,9,1,3,4,1,4,1,0,0,3,0,2,1,0,3,3,1,3,5,1,4,2,1,2,4,1,3,7,1,4,2,200,1,4,206,0,1,208,0,1,
/* out0518_em-eta18-phi25*/	13,0,2,1,0,3,2,1,3,7,1,4,2,0,0,3,0,0,1,0,3,8,0,2,1,0,3,5,1,3,3,1,4,1,200,1,2,206,0,6,
/* out0519_em-eta19-phi25*/	7,0,0,14,0,3,9,0,0,3,0,0,3,0,3,5,206,0,2,206,1,1,
/* out0520_em-eta0-phi26*/	0,
/* out0521_em-eta1-phi26*/	0,
/* out0522_em-eta2-phi26*/	0,
/* out0523_em-eta3-phi26*/	0,
/* out0524_em-eta4-phi26*/	3,12,0,4,26,1,4,26,2,1,
/* out0525_em-eta5-phi26*/	6,10,1,7,12,0,5,12,2,1,26,0,4,26,1,3,26,2,15,
/* out0526_em-eta6-phi26*/	5,8,1,2,10,0,9,10,1,1,24,1,2,24,2,12,
/* out0527_em-eta7-phi26*/	4,8,0,8,8,1,8,22,2,3,24,2,3,
/* out0528_em-eta8-phi26*/	3,6,1,9,8,0,4,22,2,5,
/* out0529_em-eta9-phi26*/	3,6,0,11,6,1,4,5,2,1,
/* out0530_em-eta10-phi26*/	9,4,1,10,6,0,2,20,2,1,5,2,15,5,3,10,5,4,7,5,5,3,5,2,8,5,5,2,
/* out0531_em-eta11-phi26*/	21,4,0,6,4,1,2,4,2,2,5,2,16,5,3,8,5,4,5,5,5,4,4,0,5,4,2,7,4,3,14,5,3,3,5,4,2,4,2,2,4,3,1,5,2,8,5,3,13,5,4,9,5,5,2,204,1,1,212,0,2,212,2,3,
/* out0532_em-eta12-phi26*/	15,2,1,5,4,0,4,4,0,2,4,2,7,4,3,14,5,3,6,5,4,4,3,2,7,4,0,7,4,0,10,4,2,5,4,3,13,204,1,8,210,2,1,212,2,5,
/* out0533_em-eta13-phi26*/	16,2,0,1,2,1,4,2,2,3,3,2,5,4,0,10,3,2,3,3,3,15,3,4,1,3,2,10,3,3,1,4,0,3,202,2,1,204,0,1,204,1,4,210,0,2,210,2,4,
/* out0534_em-eta14-phi26*/	10,2,0,4,2,2,2,3,2,5,3,3,13,2,0,2,2,3,13,2,3,5,3,3,14,202,1,8,210,0,1,
/* out0535_em-eta15-phi26*/	12,0,1,3,0,2,1,2,0,1,2,0,1,2,3,13,3,3,2,2,0,1,2,0,3,2,3,8,202,0,1,202,1,6,208,2,1,
/* out0536_em-eta16-phi26*/	9,0,1,1,0,2,3,2,0,2,1,2,1,1,3,1,200,1,2,200,2,2,202,0,1,208,0,1,
/* out0537_em-eta17-phi26*/	8,1,2,1,0,2,3,0,3,1,1,3,5,1,2,1,1,3,2,200,1,5,200,2,1,
/* out0538_em-eta18-phi26*/	8,1,3,5,0,0,1,0,2,2,0,3,2,0,3,3,1,3,4,200,0,2,200,1,3,
/* out0539_em-eta19-phi26*/	3,0,3,3,0,3,1,200,0,2,
/* out0540_em-eta0-phi27*/	0,
/* out0541_em-eta1-phi27*/	0,
/* out0542_em-eta2-phi27*/	0,
/* out0543_em-eta3-phi27*/	0,
/* out0544_em-eta4-phi27*/	2,12,0,5,12,2,1,
/* out0545_em-eta5-phi27*/	4,10,1,7,10,2,5,12,0,2,12,2,14,
/* out0546_em-eta6-phi27*/	4,8,1,2,10,0,7,10,1,1,10,2,11,
/* out0547_em-eta7-phi27*/	3,8,0,1,8,1,4,8,2,14,
/* out0548_em-eta8-phi27*/	4,6,1,3,6,2,4,8,0,3,8,2,2,
/* out0549_em-eta9-phi27*/	2,6,0,1,6,2,11,
/* out0550_em-eta10-phi27*/	5,4,1,1,4,2,4,6,0,1,6,2,1,5,3,1,
/* out0551_em-eta11-phi27*/	5,4,2,9,4,3,2,5,3,2,5,3,3,204,2,4,
/* out0552_em-eta12-phi27*/	9,2,2,1,4,0,1,4,2,1,4,3,2,5,3,2,4,3,2,204,0,2,204,1,3,204,2,8,
/* out0553_em-eta13-phi27*/	3,2,2,6,202,2,2,204,0,9,
/* out0554_em-eta14-phi27*/	3,2,2,4,202,1,1,202,2,9,
/* out0555_em-eta15-phi27*/	3,0,2,1,202,0,7,202,1,1,
/* out0556_em-eta16-phi27*/	3,0,2,3,200,2,4,202,0,3,
/* out0557_em-eta17-phi27*/	3,0,2,3,200,0,1,200,2,5,
/* out0558_em-eta18-phi27*/	1,200,0,5,
/* out0559_em-eta19-phi27*/	1,200,0,2,
/* out0560_em-eta0-phi28*/	0,
/* out0561_em-eta1-phi28*/	0,
/* out0562_em-eta2-phi28*/	0,
/* out0563_em-eta3-phi28*/	0,
/* out0564_em-eta4-phi28*/	0,
/* out0565_em-eta5-phi28*/	0,
/* out0566_em-eta6-phi28*/	0,
/* out0567_em-eta7-phi28*/	0,
/* out0568_em-eta8-phi28*/	0,
/* out0569_em-eta9-phi28*/	0,
/* out0570_em-eta10-phi28*/	0,
/* out0571_em-eta11-phi28*/	0,
/* out0572_em-eta12-phi28*/	2,204,0,2,204,2,4,
/* out0573_em-eta13-phi28*/	1,204,0,2,
/* out0574_em-eta14-phi28*/	1,202,2,4,
/* out0575_em-eta15-phi28*/	1,202,0,4,
/* out0576_em-eta16-phi28*/	1,200,2,1,
/* out0577_em-eta17-phi28*/	2,200,0,1,200,2,3,
/* out0578_em-eta18-phi28*/	1,200,0,3,
/* out0579_em-eta19-phi28*/	0,
/* out0580_em-eta0-phi29*/	0,
/* out0581_em-eta1-phi29*/	0,
/* out0582_em-eta2-phi29*/	0,
/* out0583_em-eta3-phi29*/	0,
/* out0584_em-eta4-phi29*/	0,
/* out0585_em-eta5-phi29*/	0,
/* out0586_em-eta6-phi29*/	0,
/* out0587_em-eta7-phi29*/	0,
/* out0588_em-eta8-phi29*/	0,
/* out0589_em-eta9-phi29*/	0,
/* out0590_em-eta10-phi29*/	0,
/* out0591_em-eta11-phi29*/	0,
/* out0592_em-eta12-phi29*/	0,
/* out0593_em-eta13-phi29*/	0,
/* out0594_em-eta14-phi29*/	0,
/* out0595_em-eta15-phi29*/	0,
/* out0596_em-eta16-phi29*/	0,
/* out0597_em-eta17-phi29*/	0,
/* out0598_em-eta18-phi29*/	0,
/* out0599_em-eta19-phi29*/	0
};